// vim: ts=4 sts=0 sw=0 noet
`default_nettype none
`timescale 1ns / 1ns

module ha (
	input wire [1:0] x,
	output wire [1:0] y
);
	assign y = {x[0]&x[1], x[0]^x[1]};
endmodule

module fa (
	input wire [2:0] x,
	output wire [1:0] y
);
	assign y = {(x[0]&x[1])|((x[0]^x[1])&x[2]), (x[0]^x[1])^x[2]};
endmodule

module multiplier16b (
	input wire [15:0] x, y,
	output wire [31:0] z
);
	wire [15:0][15:0] l1;

	assign l1[0] = y[0] == 0 ? '0 : x;
	assign l1[1] = y[1] == 0 ? '0 : x;
	assign l1[2] = y[2] == 0 ? '0 : x;
	assign l1[3] = y[3] == 0 ? '0 : x;
	assign l1[4] = y[4] == 0 ? '0 : x;
	assign l1[5] = y[5] == 0 ? '0 : x;
	assign l1[6] = y[6] == 0 ? '0 : x;
	assign l1[7] = y[7] == 0 ? '0 : x;
	assign l1[8] = y[8] == 0 ? '0 : x;
	assign l1[9] = y[9] == 0 ? '0 : x;
	assign l1[10] = y[10] == 0 ? '0 : x;
	assign l1[11] = y[11] == 0 ? '0 : x;
	assign l1[12] = y[12] == 0 ? '0 : x;
	assign l1[13] = y[13] == 0 ? '0 : x;
	assign l1[14] = y[14] == 0 ? '0 : x;
	assign l1[15] = y[15] == 0 ? '0 : x;

	wire l2p0 = l1[0][0];
	wire l2p1;
	wire [1:0] l2p2;
	wire [1:0] l2p3;
	wire [1:0] l2p4;
	wire [2:0] l2p5;
	wire [2:0] l2p6;
	wire [3:0] l2p7;
	wire [4:0] l2p8;
	wire [3:0] l2p9;
	wire [4:0] l2p10;
	wire [4:0] l2p11;
	wire [5:0] l2p12;
	wire [5:0] l2p13;
	wire [6:0] l2p14;
	wire [6:0] l2p15;
	wire [6:0] l2p16;
	wire [6:0] l2p17;
	wire [5:0] l2p18;
	wire [5:0] l2p19;
	wire [5:0] l2p20;
	wire [5:0] l2p21;
	wire [6:0] l2p22;
	wire [3:0] l2p23;
	wire [2:0] l2p24;
	wire [2:0] l2p25;
	wire [2:0] l2p26;
	wire [2:0] l2p27;
	wire [2:0] l2p28;
	wire [2:0] l2p29;
	wire [1:0] l2p30;

	ha hal1p1 (.x ({l1[0][1], l1[1][0]}), .y ({l2p2[0], l2p1})); // R: l2p2[0:0], l2p1
	fa fal1p2 (.x ({l1[0][2], l1[1][1], l1[2][0]}), .y ({l2p3[0], l2p2[1]})); // R: l2p3[0], l2p2[1:0]
	counter7b3 cnt7bl1p3 (
		.x ({l1[0][3], l1[1][2], l1[2][1], l1[3][0], 3'b000}),
		.y ({l2p5[0], l2p4[0], l2p3[1]})
	); // R: l2p5[0], l2p4[0], l2p3[1:0]
	counter7b3 cnt7bl1p4 (
		.x ({l1[0][4], l1[1][3], l1[2][2], l1[3][1], l1[4][0], 2'b00}),
		.y ({l2p6[0], l2p5[1], l2p4[1]})
	); // R:l2p6[0], l2p5[1:0], l2p4[1:0]
	counter7b3 cnt7bl1p5 (
		.x ({l1[0][5], l1[1][4], l1[2][3], l1[3][2], l1[4][1], l1[5][0], 1'b0}),
		.y ({l2p7[0], l2p6[1], l2p5[2]})
	); // R: l2p7[0], l2p6[1:0], l2p5[2:0]
	counter7b3 cnt7bl1p6 (
		.x ({l1[0][6], l1[1][5], l1[2][4], l1[3][3], l1[4][2], l1[5][1], l1[6][0]}),
		.y ({l2p8[0], l2p7[1], l2p6[2]})
	); // R:l2p8[0], l2p7[1:0], l2p6[2:0]
	counter7b3 cnt7bl1p7 (
		.x ({l1[0][7], l1[1][6], l1[2][5], l1[3][4], l1[4][3], l1[5][2], l1[6][1]}),
		.y ({l2p9[0], l2p8[1], l2p7[2]})
	); // R: l2p9[0], l2p8[1:0], l2p7[2:0]
	assign l2p7[3] = l1[7][0]; // R: l2p7[3:0]
	counter7b3 cnt7bl1p8 (
		.x ({l1[0][8], l1[1][7], l1[2][6], l1[3][5], l1[4][4], l1[5][3], l1[6][2]}),
		.y ({l2p10[0], l2p9[1], l2p8[2]})
	); // R: l2p10[0], l2p9[1:0], l2p8[2:0]
	assign l2p8[4:3] = {l1[7][1], l1[8][0]};
	counter7b3 cnt7bl1p9 (
		.x ({l1[0][9], l1[1][8], l1[2][7], l1[3][6], l1[4][5], l1[5][4], l1[6][3]}),
		.y ({l2p11[0], l2p10[1], l2p9[2]})
	); // R: l2p11[0], l2p10[1:0], l2p9[2:0]
	fa fal1p9 (
		.x ({l1[7][2], l1[8][1], l1[9][0]}),
		.y ({l2p10[2], l2p9[3]})
	); // R: l2p10[2:0], l2p9[3:0]
	counter7b3 cnt7bl1p10_0 (
		.x ({l1[0][10], l1[1][9], l1[2][8], l1[3][7], l1[4][6], l1[5][5], l1[6][4]}),
		.y ({l2p12[0], l2p11[1], l2p10[3]})
	); // R: l2p12[0], l2p11[1:0], l2p10[3:0]
	counter7b3 cnt7bl1p10_1 (
		.x ({l1[7][3], l1[8][2], l1[9][1], l1[10][0], 3'b000}),
		.y ({l2p12[1], l2p11[2], l2p10[4]})
	); // R: l2p12[1:0], l2p11[2:0], l2p10[4:0]
	counter7b3 cnt7bl1p11_0 (
		.x ({l1[0][11], l1[1][10], l1[2][9], l1[3][8], l1[4][7], l1[5][6], l1[6][5]}),
		.y ({l2p13[0], l2p12[2], l2p11[3]})
	); // R: l2p13[0], l2p12[2:0], l2p11[3:0]
	counter7b3 cnt7bl1p11_1 (
		.x ({l1[7][4], l1[8][3], l1[9][2], l1[10][1], l1[11][0], 2'b00}),
		.y ({l2p13[1], l2p12[3], l2p11[4]})
	); // R: l2p13[1:0], l2p12[3:0], l2p11[4:0]
	counter7b3 cnt7bl1p12_0 (
		.x ({l1[0][12], l1[1][11], l1[2][10], l1[3][9], l1[4][8], l1[5][7], l1[6][6]}),
		.y ({l2p14[0], l2p11[2], l2p12[4]})
	); // R: l2p14[0], l2p13[2:0], l2p12[4:0]
	counter7b3 cnt7bl1p12_1 (
		.x ({l1[7][5], l1[8][4], l1[9][3], l1[10][2], l1[11][1], l1[12][0], 1'b0}),
		.y ({l2p14[1], l2p13[3], l2p12[5]})
	); // R: l2p14[1:0], l2p13[3:0], l2p12[5:0]
	counter7b3 cnt7bl1p13_0 (
		.x ({l1[0][13], l1[1][12], l1[2][11], l1[3][10], l1[4][9], l1[5][8], l1[6][7]}),
		.y ({l2p15[0], l2p14[2], l2p13[4]})
	); // R: l2p15[0], l2p14[2:0], l2p13[4:0]
	counter7b3 cnt7bl1p13_1 (
		.x ({l1[7][6], l1[8][5], l1[9][4], l1[10][3], l1[11][2], l1[12][1], l1[13][0]}),
		.y ({l2p15[1], l2p14[3], l2p13[5]})
	); // R: l2p15[1:0], l2p14[3:0], l2p13[5:0]
	counter7b3 cnt7bl1p14_0 (
		.x ({l1[0][14], l1[1][13], l1[2][12], l1[3][11], l1[4][10], l1[5][9], l1[6][8]}),
		.y ({l2p16[0], l2p15[2], l2p14[4]})
	); // R: l2p16[0], l2p15[2:0], l2p14[4:0]
	counter7b3 cnt7bl1p14_1 (
		.x ({l1[7][7], l1[8][6], l1[9][5], l1[10][4], l1[11][3], l1[12][2], l1[13][1]}),
		.y ({l2p16[1], l2p15[3], l2p14[5]})
	); // R: l2p16[1:0], l2p15[3:0], l2p14[5:0]
	assign l2p14[6] = l1[14][0];
	counter7b3 cnt7bl1p15_0 (
		.x ({l1[0][15], l1[1][14], l1[2][13], l1[3][12], l1[4][11], l1[5][10], l1[6][9]}),
		.y ({l2p17[0], l2p16[2], l2p15[4]})
	); // R: l2p17[0], l2p16[2:0], l2p15[4:0]
	counter7b3 cnt7bl1p15_1 (
		.x ({l1[7][8], l1[8][7], l1[9][6], l1[10][5], l1[11][4], l1[12][3], l1[13][2]}),
		.y ({l2p17[1], l2p16[3], l2p15[5]})
	); // R: l2p17[1:0], l2p16[3:0], l2p15[5:0]


	//assign z[15:0] = x;
	//assign z[31:16] = y;
endmodule
