// vim: ts=4 sts=0 sw=0 noet
`default_nettype none
`timescale 1ns / 1ns

module testmul_tb;
	reg [15:0] x [999:0];
	reg [15:0] y [999:0];
	reg [15:0] xin;
	reg [15:0] yin;
	reg [31:0] zmul;
	wire [31:0] z;
	integer i;

	multiplier16b mul16b (
		.x (xin),
		.y (yin),
		.z (z)
	);

	initial begin
		$dumpfile("testmul_tb.vcd");
		$dumpvars(0, testmul_tb);
	end

	assign x[0] = 16'hc53e; assign y[0] = 16'hd755;
	assign x[1] = 16'h14ba; assign y[1] = 16'h8490;
	assign x[2] = 16'hf8cb; assign y[2] = 16'hcf53;
	assign x[3] = 16'h9b4b; assign y[3] = 16'hf404;
	assign x[4] = 16'hb752; assign y[4] = 16'h6fd7;
	assign x[5] = 16'h474e; assign y[5] = 16'h904d;
	assign x[6] = 16'h478c; assign y[6] = 16'h308d;
	assign x[7] = 16'h8042; assign y[7] = 16'h4b3e;
	assign x[8] = 16'h9ecb; assign y[8] = 16'h3291;
	assign x[9] = 16'h25c1; assign y[9] = 16'ha90f;
	assign x[10] = 16'hf1bc; assign y[10] = 16'h338f;
	assign x[11] = 16'hb524; assign y[11] = 16'hde4b;
	assign x[12] = 16'ha1e4; assign y[12] = 16'h68b1;
	assign x[13] = 16'hf43a; assign y[13] = 16'he2a8;
	assign x[14] = 16'h855f; assign y[14] = 16'h1fe3;
	assign x[15] = 16'h0730; assign y[15] = 16'h2fc1;
	assign x[16] = 16'hcc32; assign y[16] = 16'h0095;
	assign x[17] = 16'hfcb6; assign y[17] = 16'haa90;
	assign x[18] = 16'h7ce1; assign y[18] = 16'ha681;
	assign x[19] = 16'h203f; assign y[19] = 16'h61d3;
	assign x[20] = 16'h7183; assign y[20] = 16'h7a2b;
	assign x[21] = 16'h48f5; assign y[21] = 16'he55c;
	assign x[22] = 16'h2eb3; assign y[22] = 16'h2930;
	assign x[23] = 16'ha3de; assign y[23] = 16'hfa83;
	assign x[24] = 16'h37d6; assign y[24] = 16'h9a57;
	assign x[25] = 16'h9509; assign y[25] = 16'h3fe7;
	assign x[26] = 16'haa5e; assign y[26] = 16'h680a;
	assign x[27] = 16'h9347; assign y[27] = 16'he3d5;
	assign x[28] = 16'h2eea; assign y[28] = 16'hc511;
	assign x[29] = 16'ha253; assign y[29] = 16'h7bf5;
	assign x[30] = 16'h94a6; assign y[30] = 16'h5e24;
	assign x[31] = 16'h60f7; assign y[31] = 16'h5f9b;
	assign x[32] = 16'h10e1; assign y[32] = 16'h8526;
	assign x[33] = 16'hf3fb; assign y[33] = 16'h235f;
	assign x[34] = 16'h2dfd; assign y[34] = 16'h42ac;
	assign x[35] = 16'h4c91; assign y[35] = 16'h13c8;
	assign x[36] = 16'h2916; assign y[36] = 16'hc857;
	assign x[37] = 16'h8d1f; assign y[37] = 16'h7893;
	assign x[38] = 16'h6e2e; assign y[38] = 16'hd6be;
	assign x[39] = 16'h8ce8; assign y[39] = 16'he6b0;
	assign x[40] = 16'hfc3d; assign y[40] = 16'hb6f8;
	assign x[41] = 16'h2a2c; assign y[41] = 16'ha60d;
	assign x[42] = 16'h3b0f; assign y[42] = 16'hf90f;
	assign x[43] = 16'haba8; assign y[43] = 16'h6179;
	assign x[44] = 16'h7c6f; assign y[44] = 16'h084c;
	assign x[45] = 16'h8ac5; assign y[45] = 16'h3bf9;
	assign x[46] = 16'h70e0; assign y[46] = 16'hbe7e;
	assign x[47] = 16'h5749; assign y[47] = 16'haa42;
	assign x[48] = 16'hda2d; assign y[48] = 16'h1fd7;
	assign x[49] = 16'h3382; assign y[49] = 16'h4aef;
	assign x[50] = 16'h7003; assign y[50] = 16'h1728;
	assign x[51] = 16'h25e2; assign y[51] = 16'h0dab;
	assign x[52] = 16'h3fb7; assign y[52] = 16'h6085;
	assign x[53] = 16'h3d48; assign y[53] = 16'hc84c;
	assign x[54] = 16'h2edd; assign y[54] = 16'hbd82;
	assign x[55] = 16'h3b6a; assign y[55] = 16'h12a1;
	assign x[56] = 16'h0b13; assign y[56] = 16'h63a1;
	assign x[57] = 16'h5eb4; assign y[57] = 16'h3f6f;
	assign x[58] = 16'hf55e; assign y[58] = 16'h6bd0;
	assign x[59] = 16'h1f46; assign y[59] = 16'h0baa;
	assign x[60] = 16'hd9ea; assign y[60] = 16'h33f7;
	assign x[61] = 16'h8514; assign y[61] = 16'h23d7;
	assign x[62] = 16'h7110; assign y[62] = 16'h24d9;
	assign x[63] = 16'h9a24; assign y[63] = 16'hb359;
	assign x[64] = 16'hdf44; assign y[64] = 16'h5c52;
	assign x[65] = 16'h1f40; assign y[65] = 16'hef2b;
	assign x[66] = 16'h1429; assign y[66] = 16'h33ab;
	assign x[67] = 16'hc855; assign y[67] = 16'h6611;
	assign x[68] = 16'h8530; assign y[68] = 16'hb794;
	assign x[69] = 16'hf0c0; assign y[69] = 16'h56be;
	assign x[70] = 16'h6825; assign y[70] = 16'h1db8;
	assign x[71] = 16'h5100; assign y[71] = 16'h52eb;
	assign x[72] = 16'haf43; assign y[72] = 16'h805a;
	assign x[73] = 16'h3c03; assign y[73] = 16'he276;
	assign x[74] = 16'h5981; assign y[74] = 16'h06c2;
	assign x[75] = 16'hf178; assign y[75] = 16'hd1df;
	assign x[76] = 16'h9f75; assign y[76] = 16'hb6dc;
	assign x[77] = 16'hc6fc; assign y[77] = 16'h807a;
	assign x[78] = 16'h4e8c; assign y[78] = 16'h065e;
	assign x[79] = 16'hea78; assign y[79] = 16'h287c;
	assign x[80] = 16'habfd; assign y[80] = 16'h1765;
	assign x[81] = 16'h8fcf; assign y[81] = 16'h4509;
	assign x[82] = 16'h7af2; assign y[82] = 16'hf6b2;
	assign x[83] = 16'hb456; assign y[83] = 16'h9364;
	assign x[84] = 16'hb7e9; assign y[84] = 16'h43c2;
	assign x[85] = 16'h9edf; assign y[85] = 16'hc6aa;
	assign x[86] = 16'hd42e; assign y[86] = 16'h2954;
	assign x[87] = 16'h00c7; assign y[87] = 16'h6276;
	assign x[88] = 16'hab36; assign y[88] = 16'h51f5;
	assign x[89] = 16'h7a94; assign y[89] = 16'h7239;
	assign x[90] = 16'he571; assign y[90] = 16'hc1de;
	assign x[91] = 16'hd42d; assign y[91] = 16'h1026;
	assign x[92] = 16'hcdf5; assign y[92] = 16'hd621;
	assign x[93] = 16'h17f3; assign y[93] = 16'h54d3;
	assign x[94] = 16'he405; assign y[94] = 16'h20b5;
	assign x[95] = 16'h84b9; assign y[95] = 16'h50bc;
	assign x[96] = 16'he489; assign y[96] = 16'hf97a;
	assign x[97] = 16'h0009; assign y[97] = 16'h13ec;
	assign x[98] = 16'hfd39; assign y[98] = 16'ha6e2;
	assign x[99] = 16'h9fc6; assign y[99] = 16'hef0c;
	assign x[100] = 16'h1986; assign y[100] = 16'hd48c;
	assign x[101] = 16'h6041; assign y[101] = 16'h2abc;
	assign x[102] = 16'h42d3; assign y[102] = 16'h078a;
	assign x[103] = 16'hcdba; assign y[103] = 16'hd5c0;
	assign x[104] = 16'ha1e1; assign y[104] = 16'h01bc;
	assign x[105] = 16'h6d53; assign y[105] = 16'h0751;
	assign x[106] = 16'h0135; assign y[106] = 16'h3210;
	assign x[107] = 16'h6183; assign y[107] = 16'h3ce0;
	assign x[108] = 16'h65a3; assign y[108] = 16'h9ad6;
	assign x[109] = 16'h8f59; assign y[109] = 16'h5d4c;
	assign x[110] = 16'h334a; assign y[110] = 16'hf382;
	assign x[111] = 16'hcb1b; assign y[111] = 16'h29a6;
	assign x[112] = 16'h0b2f; assign y[112] = 16'h8ca7;
	assign x[113] = 16'he7ec; assign y[113] = 16'h3b47;
	assign x[114] = 16'h8352; assign y[114] = 16'h444f;
	assign x[115] = 16'hb1b0; assign y[115] = 16'h3aef;
	assign x[116] = 16'h4f12; assign y[116] = 16'h8e8b;
	assign x[117] = 16'h0982; assign y[117] = 16'h15a8;
	assign x[118] = 16'h14d1; assign y[118] = 16'h6956;
	assign x[119] = 16'h84f3; assign y[119] = 16'ha122;
	assign x[120] = 16'hbbd9; assign y[120] = 16'h1581;
	assign x[121] = 16'hfd2d; assign y[121] = 16'head6;
	assign x[122] = 16'hdef2; assign y[122] = 16'hbeb1;
	assign x[123] = 16'h5b48; assign y[123] = 16'h6a6a;
	assign x[124] = 16'hc04b; assign y[124] = 16'h9502;
	assign x[125] = 16'h048e; assign y[125] = 16'h46e3;
	assign x[126] = 16'h4d52; assign y[126] = 16'h8af1;
	assign x[127] = 16'haab4; assign y[127] = 16'hacce;
	assign x[128] = 16'hbc01; assign y[128] = 16'h2ffa;
	assign x[129] = 16'had2f; assign y[129] = 16'h1242;
	assign x[130] = 16'h1518; assign y[130] = 16'h8a0b;
	assign x[131] = 16'h53e5; assign y[131] = 16'h4c80;
	assign x[132] = 16'h943d; assign y[132] = 16'hb8c8;
	assign x[133] = 16'hca22; assign y[133] = 16'h4260;
	assign x[134] = 16'h9639; assign y[134] = 16'h3ad3;
	assign x[135] = 16'hf4c4; assign y[135] = 16'h7aba;
	assign x[136] = 16'h18b5; assign y[136] = 16'h9da2;
	assign x[137] = 16'h5bf2; assign y[137] = 16'h2448;
	assign x[138] = 16'h9af7; assign y[138] = 16'hce6c;
	assign x[139] = 16'ha833; assign y[139] = 16'h9934;
	assign x[140] = 16'hd456; assign y[140] = 16'h37a1;
	assign x[141] = 16'h32e4; assign y[141] = 16'hf65c;
	assign x[142] = 16'hf2b0; assign y[142] = 16'hac95;
	assign x[143] = 16'haff3; assign y[143] = 16'h3fa7;
	assign x[144] = 16'hf54a; assign y[144] = 16'h3b65;
	assign x[145] = 16'hfed7; assign y[145] = 16'hda62;
	assign x[146] = 16'h135d; assign y[146] = 16'h9a93;
	assign x[147] = 16'hab8f; assign y[147] = 16'h4fb3;
	assign x[148] = 16'h5546; assign y[148] = 16'hc04a;
	assign x[149] = 16'h2c81; assign y[149] = 16'h21b5;
	assign x[150] = 16'h2b59; assign y[150] = 16'h6565;
	assign x[151] = 16'h712e; assign y[151] = 16'h1f4f;
	assign x[152] = 16'hc506; assign y[152] = 16'h0405;
	assign x[153] = 16'h3237; assign y[153] = 16'hc9a1;
	assign x[154] = 16'h9463; assign y[154] = 16'he5a7;
	assign x[155] = 16'hfa2c; assign y[155] = 16'h6f3b;
	assign x[156] = 16'hd898; assign y[156] = 16'h2ad5;
	assign x[157] = 16'hbc95; assign y[157] = 16'h70b5;
	assign x[158] = 16'h8596; assign y[158] = 16'h554a;
	assign x[159] = 16'hdcc9; assign y[159] = 16'h6246;
	assign x[160] = 16'hb78f; assign y[160] = 16'h3ae2;
	assign x[161] = 16'h20b1; assign y[161] = 16'h0e24;
	assign x[162] = 16'he739; assign y[162] = 16'h6743;
	assign x[163] = 16'h3ce1; assign y[163] = 16'hfe82;
	assign x[164] = 16'hcbc0; assign y[164] = 16'h8351;
	assign x[165] = 16'h6a1a; assign y[165] = 16'h158e;
	assign x[166] = 16'h6e89; assign y[166] = 16'h4aee;
	assign x[167] = 16'h3592; assign y[167] = 16'h655c;
	assign x[168] = 16'heab4; assign y[168] = 16'hc18d;
	assign x[169] = 16'hb929; assign y[169] = 16'h4d7b;
	assign x[170] = 16'h35a1; assign y[170] = 16'hf9ce;
	assign x[171] = 16'h4bfb; assign y[171] = 16'hcfd3;
	assign x[172] = 16'hd8b2; assign y[172] = 16'hfda5;
	assign x[173] = 16'ha519; assign y[173] = 16'hff33;
	assign x[174] = 16'hff4e; assign y[174] = 16'h676b;
	assign x[175] = 16'h7003; assign y[175] = 16'h04f8;
	assign x[176] = 16'hae31; assign y[176] = 16'ha2f2;
	assign x[177] = 16'ha4c6; assign y[177] = 16'h1228;
	assign x[178] = 16'h4bf6; assign y[178] = 16'h8386;
	assign x[179] = 16'h4fd2; assign y[179] = 16'hc20c;
	assign x[180] = 16'h96b9; assign y[180] = 16'hf0dc;
	assign x[181] = 16'h21f9; assign y[181] = 16'h2b56;
	assign x[182] = 16'h142e; assign y[182] = 16'h21f9;
	assign x[183] = 16'h733f; assign y[183] = 16'h42d0;
	assign x[184] = 16'h14cd; assign y[184] = 16'h99d4;
	assign x[185] = 16'h07d3; assign y[185] = 16'he5ad;
	assign x[186] = 16'ha943; assign y[186] = 16'h5245;
	assign x[187] = 16'h4c32; assign y[187] = 16'hebe5;
	assign x[188] = 16'hbe1d; assign y[188] = 16'hc3b3;
	assign x[189] = 16'h1136; assign y[189] = 16'h2e69;
	assign x[190] = 16'h2718; assign y[190] = 16'hda4c;
	assign x[191] = 16'h6986; assign y[191] = 16'h944e;
	assign x[192] = 16'hd5ef; assign y[192] = 16'hf6e4;
	assign x[193] = 16'hc6f2; assign y[193] = 16'h7796;
	assign x[194] = 16'h0a7c; assign y[194] = 16'h001f;
	assign x[195] = 16'h5d2b; assign y[195] = 16'h9ad9;
	assign x[196] = 16'h8248; assign y[196] = 16'haa55;
	assign x[197] = 16'h2199; assign y[197] = 16'hfcad;
	assign x[198] = 16'h8625; assign y[198] = 16'h9b09;
	assign x[199] = 16'hd0ee; assign y[199] = 16'hc4b0;
	assign x[200] = 16'hc471; assign y[200] = 16'h1fe0;
	assign x[201] = 16'h53dc; assign y[201] = 16'h4130;
	assign x[202] = 16'h7a57; assign y[202] = 16'h92fd;
	assign x[203] = 16'hab05; assign y[203] = 16'h1c6e;
	assign x[204] = 16'h1265; assign y[204] = 16'hf670;
	assign x[205] = 16'hd5f2; assign y[205] = 16'h4824;
	assign x[206] = 16'hfbd1; assign y[206] = 16'h29ca;
	assign x[207] = 16'h4d80; assign y[207] = 16'hb49e;
	assign x[208] = 16'hd280; assign y[208] = 16'h1203;
	assign x[209] = 16'heebc; assign y[209] = 16'hc5fb;
	assign x[210] = 16'heaf2; assign y[210] = 16'h1814;
	assign x[211] = 16'h33f5; assign y[211] = 16'hf118;
	assign x[212] = 16'h4d80; assign y[212] = 16'h0a5b;
	assign x[213] = 16'h109f; assign y[213] = 16'h43f1;
	assign x[214] = 16'ha5d7; assign y[214] = 16'h35e8;
	assign x[215] = 16'hb17e; assign y[215] = 16'h63d3;
	assign x[216] = 16'hc44e; assign y[216] = 16'hfb0b;
	assign x[217] = 16'h38d4; assign y[217] = 16'h1ecd;
	assign x[218] = 16'hef33; assign y[218] = 16'hacfc;
	assign x[219] = 16'h3fa7; assign y[219] = 16'h97bf;
	assign x[220] = 16'h4114; assign y[220] = 16'hc679;
	assign x[221] = 16'h966d; assign y[221] = 16'h3e3c;
	assign x[222] = 16'h60d5; assign y[222] = 16'h138c;
	assign x[223] = 16'hc8b7; assign y[223] = 16'he39f;
	assign x[224] = 16'hbe3f; assign y[224] = 16'h6186;
	assign x[225] = 16'he933; assign y[225] = 16'hb68e;
	assign x[226] = 16'h2692; assign y[226] = 16'h16db;
	assign x[227] = 16'h1478; assign y[227] = 16'hf8ea;
	assign x[228] = 16'h82c1; assign y[228] = 16'h0da5;
	assign x[229] = 16'h6e94; assign y[229] = 16'h7595;
	assign x[230] = 16'h2fdc; assign y[230] = 16'hd718;
	assign x[231] = 16'h9c51; assign y[231] = 16'h3a15;
	assign x[232] = 16'h4a97; assign y[232] = 16'hda18;
	assign x[233] = 16'hd817; assign y[233] = 16'h2b06;
	assign x[234] = 16'h35a3; assign y[234] = 16'hd4ce;
	assign x[235] = 16'h2037; assign y[235] = 16'h32cb;
	assign x[236] = 16'hd490; assign y[236] = 16'h4ff3;
	assign x[237] = 16'h0fb8; assign y[237] = 16'he4b8;
	assign x[238] = 16'hdcb7; assign y[238] = 16'hd583;
	assign x[239] = 16'h0f6d; assign y[239] = 16'hfe45;
	assign x[240] = 16'ha624; assign y[240] = 16'h8152;
	assign x[241] = 16'h2836; assign y[241] = 16'hb47b;
	assign x[242] = 16'h2402; assign y[242] = 16'h3e25;
	assign x[243] = 16'hb7f0; assign y[243] = 16'h0f0a;
	assign x[244] = 16'hb0de; assign y[244] = 16'hb21d;
	assign x[245] = 16'h5b16; assign y[245] = 16'h051a;
	assign x[246] = 16'h7603; assign y[246] = 16'hbb4a;
	assign x[247] = 16'h241a; assign y[247] = 16'h495d;
	assign x[248] = 16'h6a7c; assign y[248] = 16'h01a7;
	assign x[249] = 16'h68da; assign y[249] = 16'h3f12;
	assign x[250] = 16'h03ad; assign y[250] = 16'h9626;
	assign x[251] = 16'hbcfe; assign y[251] = 16'h0c9e;
	assign x[252] = 16'h7739; assign y[252] = 16'h48a5;
	assign x[253] = 16'h5fbd; assign y[253] = 16'he878;
	assign x[254] = 16'h398b; assign y[254] = 16'hf411;
	assign x[255] = 16'hb05b; assign y[255] = 16'h8435;
	assign x[256] = 16'h42a4; assign y[256] = 16'h0e4d;
	assign x[257] = 16'h6a8e; assign y[257] = 16'hb977;
	assign x[258] = 16'hab86; assign y[258] = 16'hf25d;
	assign x[259] = 16'h95d3; assign y[259] = 16'h97ba;
	assign x[260] = 16'ha76a; assign y[260] = 16'h5e3b;
	assign x[261] = 16'h295f; assign y[261] = 16'h3485;
	assign x[262] = 16'h9d93; assign y[262] = 16'h5014;
	assign x[263] = 16'hc0d0; assign y[263] = 16'h4b39;
	assign x[264] = 16'h401e; assign y[264] = 16'h7215;
	assign x[265] = 16'ha1bc; assign y[265] = 16'h7c55;
	assign x[266] = 16'h792b; assign y[266] = 16'h5e2d;
	assign x[267] = 16'h9505; assign y[267] = 16'hbeb3;
	assign x[268] = 16'hd6ee; assign y[268] = 16'h17ae;
	assign x[269] = 16'h43b4; assign y[269] = 16'h0a85;
	assign x[270] = 16'hc9a0; assign y[270] = 16'h27e5;
	assign x[271] = 16'h257b; assign y[271] = 16'h4398;
	assign x[272] = 16'hd728; assign y[272] = 16'h9949;
	assign x[273] = 16'hd560; assign y[273] = 16'h48d9;
	assign x[274] = 16'hd829; assign y[274] = 16'h9897;
	assign x[275] = 16'hb589; assign y[275] = 16'h2b4a;
	assign x[276] = 16'h7f01; assign y[276] = 16'he3be;
	assign x[277] = 16'hbd0f; assign y[277] = 16'h1d9f;
	assign x[278] = 16'hc0bb; assign y[278] = 16'hd137;
	assign x[279] = 16'h0450; assign y[279] = 16'hd59e;
	assign x[280] = 16'ha42e; assign y[280] = 16'he1f1;
	assign x[281] = 16'h6871; assign y[281] = 16'hbe41;
	assign x[282] = 16'h962c; assign y[282] = 16'hf118;
	assign x[283] = 16'h2e9e; assign y[283] = 16'h5ef4;
	assign x[284] = 16'h379c; assign y[284] = 16'h8dcf;
	assign x[285] = 16'h396c; assign y[285] = 16'h4ec9;
	assign x[286] = 16'he46f; assign y[286] = 16'hcc2c;
	assign x[287] = 16'h5eea; assign y[287] = 16'hd7e9;
	assign x[288] = 16'hdd09; assign y[288] = 16'h5977;
	assign x[289] = 16'h7ef4; assign y[289] = 16'he82a;
	assign x[290] = 16'hae47; assign y[290] = 16'h48fe;
	assign x[291] = 16'hb5f2; assign y[291] = 16'hecc4;
	assign x[292] = 16'h2c49; assign y[292] = 16'hf771;
	assign x[293] = 16'h6843; assign y[293] = 16'h96e6;
	assign x[294] = 16'h00f1; assign y[294] = 16'he5ee;
	assign x[295] = 16'hec8c; assign y[295] = 16'h03fb;
	assign x[296] = 16'h6ffd; assign y[296] = 16'h98dc;
	assign x[297] = 16'h3a9a; assign y[297] = 16'h9a31;
	assign x[298] = 16'h4ffc; assign y[298] = 16'hd931;
	assign x[299] = 16'hf15f; assign y[299] = 16'h2f63;
	assign x[300] = 16'hfecf; assign y[300] = 16'h76f8;
	assign x[301] = 16'hcf84; assign y[301] = 16'h8f67;
	assign x[302] = 16'h0b11; assign y[302] = 16'h3ddd;
	assign x[303] = 16'h8a47; assign y[303] = 16'h14c2;
	assign x[304] = 16'h0021; assign y[304] = 16'h835d;
	assign x[305] = 16'hcbfe; assign y[305] = 16'hcadf;
	assign x[306] = 16'he3a0; assign y[306] = 16'h343d;
	assign x[307] = 16'h8155; assign y[307] = 16'hb528;
	assign x[308] = 16'h9119; assign y[308] = 16'h645e;
	assign x[309] = 16'h2ba7; assign y[309] = 16'h1226;
	assign x[310] = 16'h2412; assign y[310] = 16'h8664;
	assign x[311] = 16'h9c78; assign y[311] = 16'hae06;
	assign x[312] = 16'h3c82; assign y[312] = 16'h7f83;
	assign x[313] = 16'h53bd; assign y[313] = 16'h22dd;
	assign x[314] = 16'hd464; assign y[314] = 16'h9452;
	assign x[315] = 16'h90c4; assign y[315] = 16'h44d2;
	assign x[316] = 16'h6ba9; assign y[316] = 16'h35ea;
	assign x[317] = 16'hd254; assign y[317] = 16'hce8c;
	assign x[318] = 16'h8ea6; assign y[318] = 16'h95a2;
	assign x[319] = 16'he27d; assign y[319] = 16'hbe5d;
	assign x[320] = 16'h468f; assign y[320] = 16'h506b;
	assign x[321] = 16'h3f20; assign y[321] = 16'h3db4;
	assign x[322] = 16'hc34a; assign y[322] = 16'hcd6c;
	assign x[323] = 16'hef96; assign y[323] = 16'h4770;
	assign x[324] = 16'h9911; assign y[324] = 16'hb547;
	assign x[325] = 16'hf201; assign y[325] = 16'hd488;
	assign x[326] = 16'h6f9f; assign y[326] = 16'hf414;
	assign x[327] = 16'hfa4b; assign y[327] = 16'ha2f0;
	assign x[328] = 16'hfc45; assign y[328] = 16'h1ed5;
	assign x[329] = 16'he351; assign y[329] = 16'h99b1;
	assign x[330] = 16'h491e; assign y[330] = 16'hfdb5;
	assign x[331] = 16'h1ad4; assign y[331] = 16'h6e72;
	assign x[332] = 16'h0d14; assign y[332] = 16'hb5f7;
	assign x[333] = 16'hf16c; assign y[333] = 16'hc82c;
	assign x[334] = 16'h052d; assign y[334] = 16'h2206;
	assign x[335] = 16'h29a9; assign y[335] = 16'hca4c;
	assign x[336] = 16'h0349; assign y[336] = 16'hb8f9;
	assign x[337] = 16'h1515; assign y[337] = 16'h3b78;
	assign x[338] = 16'h01ea; assign y[338] = 16'h8a68;
	assign x[339] = 16'h95c6; assign y[339] = 16'h7410;
	assign x[340] = 16'h4807; assign y[340] = 16'h936a;
	assign x[341] = 16'h61e5; assign y[341] = 16'h35fe;
	assign x[342] = 16'hde37; assign y[342] = 16'hebfa;
	assign x[343] = 16'ha90f; assign y[343] = 16'hc4ac;
	assign x[344] = 16'h5625; assign y[344] = 16'ha950;
	assign x[345] = 16'hd7ea; assign y[345] = 16'hdedb;
	assign x[346] = 16'h4bc9; assign y[346] = 16'he503;
	assign x[347] = 16'h4b85; assign y[347] = 16'ha1d4;
	assign x[348] = 16'h4229; assign y[348] = 16'h6af0;
	assign x[349] = 16'h5fa7; assign y[349] = 16'he364;
	assign x[350] = 16'hb2c6; assign y[350] = 16'hc71a;
	assign x[351] = 16'hdac5; assign y[351] = 16'hfbe1;
	assign x[352] = 16'hc771; assign y[352] = 16'h70b8;
	assign x[353] = 16'h6473; assign y[353] = 16'he0e8;
	assign x[354] = 16'h6895; assign y[354] = 16'h197e;
	assign x[355] = 16'hc6d5; assign y[355] = 16'h1109;
	assign x[356] = 16'h77d2; assign y[356] = 16'h2b58;
	assign x[357] = 16'h5f9e; assign y[357] = 16'hba2b;
	assign x[358] = 16'h1d2d; assign y[358] = 16'h58c4;
	assign x[359] = 16'h7754; assign y[359] = 16'h9855;
	assign x[360] = 16'h2c5a; assign y[360] = 16'h91a0;
	assign x[361] = 16'hb4c5; assign y[361] = 16'hd2a7;
	assign x[362] = 16'heaa5; assign y[362] = 16'h1b9e;
	assign x[363] = 16'hdc78; assign y[363] = 16'he8c1;
	assign x[364] = 16'hfafb; assign y[364] = 16'h826e;
	assign x[365] = 16'hf388; assign y[365] = 16'h6e4b;
	assign x[366] = 16'haca4; assign y[366] = 16'h8820;
	assign x[367] = 16'h159f; assign y[367] = 16'h166d;
	assign x[368] = 16'h1ae8; assign y[368] = 16'h5362;
	assign x[369] = 16'hb319; assign y[369] = 16'h01fb;
	assign x[370] = 16'h9461; assign y[370] = 16'h03a6;
	assign x[371] = 16'h47e3; assign y[371] = 16'h209b;
	assign x[372] = 16'hdb01; assign y[372] = 16'h71bf;
	assign x[373] = 16'hcb03; assign y[373] = 16'h7123;
	assign x[374] = 16'he84b; assign y[374] = 16'h62bd;
	assign x[375] = 16'hadd3; assign y[375] = 16'h3465;
	assign x[376] = 16'h2bd6; assign y[376] = 16'ha357;
	assign x[377] = 16'ha556; assign y[377] = 16'he957;
	assign x[378] = 16'ha679; assign y[378] = 16'h82d0;
	assign x[379] = 16'h0ec2; assign y[379] = 16'h16b5;
	assign x[380] = 16'h6158; assign y[380] = 16'hbcc6;
	assign x[381] = 16'h2904; assign y[381] = 16'h6b4f;
	assign x[382] = 16'hb105; assign y[382] = 16'h6025;
	assign x[383] = 16'h673a; assign y[383] = 16'h80a7;
	assign x[384] = 16'h9a46; assign y[384] = 16'h9fdc;
	assign x[385] = 16'hc4f3; assign y[385] = 16'h8260;
	assign x[386] = 16'hf6d3; assign y[386] = 16'hb018;
	assign x[387] = 16'h7adc; assign y[387] = 16'h16c9;
	assign x[388] = 16'h9c93; assign y[388] = 16'h2509;
	assign x[389] = 16'h04b6; assign y[389] = 16'hebff;
	assign x[390] = 16'hfd98; assign y[390] = 16'he05b;
	assign x[391] = 16'h184d; assign y[391] = 16'hd301;
	assign x[392] = 16'hfcb6; assign y[392] = 16'hebc8;
	assign x[393] = 16'he155; assign y[393] = 16'h3c7a;
	assign x[394] = 16'h2bd5; assign y[394] = 16'h29b7;
	assign x[395] = 16'h7b77; assign y[395] = 16'h328c;
	assign x[396] = 16'h4ebe; assign y[396] = 16'hd3f9;
	assign x[397] = 16'h6d4b; assign y[397] = 16'he19b;
	assign x[398] = 16'h277f; assign y[398] = 16'hda97;
	assign x[399] = 16'hc9f8; assign y[399] = 16'h1425;
	assign x[400] = 16'h5c5b; assign y[400] = 16'h7fdc;
	assign x[401] = 16'hfae3; assign y[401] = 16'h70aa;
	assign x[402] = 16'h4194; assign y[402] = 16'h8ed8;
	assign x[403] = 16'hb446; assign y[403] = 16'ha3a2;
	assign x[404] = 16'hdea3; assign y[404] = 16'h36ee;
	assign x[405] = 16'h922d; assign y[405] = 16'h6701;
	assign x[406] = 16'h97e1; assign y[406] = 16'he231;
	assign x[407] = 16'hec95; assign y[407] = 16'h85a0;
	assign x[408] = 16'h8b8b; assign y[408] = 16'h76ac;
	assign x[409] = 16'h087a; assign y[409] = 16'h3cca;
	assign x[410] = 16'h32a3; assign y[410] = 16'h585b;
	assign x[411] = 16'hd44e; assign y[411] = 16'h7f5f;
	assign x[412] = 16'h6fa6; assign y[412] = 16'h91b1;
	assign x[413] = 16'h034c; assign y[413] = 16'hdb46;
	assign x[414] = 16'h197b; assign y[414] = 16'h3e5b;
	assign x[415] = 16'hc4f6; assign y[415] = 16'h8b83;
	assign x[416] = 16'h3c8a; assign y[416] = 16'hb7c2;
	assign x[417] = 16'h7589; assign y[417] = 16'h9078;
	assign x[418] = 16'h7170; assign y[418] = 16'h7af3;
	assign x[419] = 16'h212b; assign y[419] = 16'h9d73;
	assign x[420] = 16'ha795; assign y[420] = 16'h779a;
	assign x[421] = 16'hbf13; assign y[421] = 16'hf5e5;
	assign x[422] = 16'h92db; assign y[422] = 16'h57bf;
	assign x[423] = 16'h464a; assign y[423] = 16'h07ef;
	assign x[424] = 16'ha7e0; assign y[424] = 16'hbbe5;
	assign x[425] = 16'h0cf2; assign y[425] = 16'h4278;
	assign x[426] = 16'hca89; assign y[426] = 16'h4f7c;
	assign x[427] = 16'h5a80; assign y[427] = 16'h2725;
	assign x[428] = 16'h456a; assign y[428] = 16'h69ba;
	assign x[429] = 16'hfe54; assign y[429] = 16'h6d4a;
	assign x[430] = 16'h787b; assign y[430] = 16'h43a6;
	assign x[431] = 16'h77a6; assign y[431] = 16'hc4eb;
	assign x[432] = 16'hb4f9; assign y[432] = 16'h43dc;
	assign x[433] = 16'hff36; assign y[433] = 16'h374d;
	assign x[434] = 16'h0d51; assign y[434] = 16'hb79c;
	assign x[435] = 16'hfa78; assign y[435] = 16'he944;
	assign x[436] = 16'h9e0d; assign y[436] = 16'h0678;
	assign x[437] = 16'h70ad; assign y[437] = 16'h5379;
	assign x[438] = 16'hfd49; assign y[438] = 16'hf63a;
	assign x[439] = 16'ha0bd; assign y[439] = 16'h2854;
	assign x[440] = 16'h84b0; assign y[440] = 16'h465f;
	assign x[441] = 16'hcdbf; assign y[441] = 16'h61d3;
	assign x[442] = 16'ha201; assign y[442] = 16'h955d;
	assign x[443] = 16'hc4a7; assign y[443] = 16'h1e4c;
	assign x[444] = 16'h6ad5; assign y[444] = 16'h139a;
	assign x[445] = 16'ha15c; assign y[445] = 16'h7fcc;
	assign x[446] = 16'hafb3; assign y[446] = 16'he1e4;
	assign x[447] = 16'h73ab; assign y[447] = 16'h852c;
	assign x[448] = 16'hb037; assign y[448] = 16'h531d;
	assign x[449] = 16'h9c1c; assign y[449] = 16'h08b1;
	assign x[450] = 16'hb674; assign y[450] = 16'h1dca;
	assign x[451] = 16'h4d6c; assign y[451] = 16'hb4f3;
	assign x[452] = 16'h0b41; assign y[452] = 16'hfb72;
	assign x[453] = 16'h1f65; assign y[453] = 16'h0c93;
	assign x[454] = 16'h7ba1; assign y[454] = 16'h1705;
	assign x[455] = 16'h065e; assign y[455] = 16'h7398;
	assign x[456] = 16'ha741; assign y[456] = 16'h2212;
	assign x[457] = 16'h1ff3; assign y[457] = 16'hb09a;
	assign x[458] = 16'hd865; assign y[458] = 16'h458e;
	assign x[459] = 16'h6edc; assign y[459] = 16'he5de;
	assign x[460] = 16'hded4; assign y[460] = 16'h48bb;
	assign x[461] = 16'hb750; assign y[461] = 16'h9fb8;
	assign x[462] = 16'h5a97; assign y[462] = 16'ha85a;
	assign x[463] = 16'hd138; assign y[463] = 16'hc3ed;
	assign x[464] = 16'h04ee; assign y[464] = 16'hd18d;
	assign x[465] = 16'h8709; assign y[465] = 16'hece0;
	assign x[466] = 16'h1579; assign y[466] = 16'h3ec4;
	assign x[467] = 16'hd15f; assign y[467] = 16'hc7d5;
	assign x[468] = 16'h57b6; assign y[468] = 16'h0197;
	assign x[469] = 16'h46c5; assign y[469] = 16'h4bdc;
	assign x[470] = 16'h28c7; assign y[470] = 16'ha8fc;
	assign x[471] = 16'h7989; assign y[471] = 16'h5a40;
	assign x[472] = 16'h7e5b; assign y[472] = 16'h0b40;
	assign x[473] = 16'h5672; assign y[473] = 16'h562d;
	assign x[474] = 16'h282f; assign y[474] = 16'hdab6;
	assign x[475] = 16'h3512; assign y[475] = 16'hea3e;
	assign x[476] = 16'h4cd6; assign y[476] = 16'h1481;
	assign x[477] = 16'h8144; assign y[477] = 16'hae35;
	assign x[478] = 16'hc0c6; assign y[478] = 16'h0df5;
	assign x[479] = 16'h1298; assign y[479] = 16'hfe20;
	assign x[480] = 16'h2de2; assign y[480] = 16'hb77b;
	assign x[481] = 16'h95e1; assign y[481] = 16'h4d36;
	assign x[482] = 16'hea8e; assign y[482] = 16'h78e8;
	assign x[483] = 16'hb62c; assign y[483] = 16'h5316;
	assign x[484] = 16'hcf36; assign y[484] = 16'hacdf;
	assign x[485] = 16'h8a28; assign y[485] = 16'hfc10;
	assign x[486] = 16'hc901; assign y[486] = 16'h0791;
	assign x[487] = 16'h9f1c; assign y[487] = 16'h9392;
	assign x[488] = 16'hf015; assign y[488] = 16'h11e2;
	assign x[489] = 16'h865f; assign y[489] = 16'h139c;
	assign x[490] = 16'he96e; assign y[490] = 16'hca45;
	assign x[491] = 16'h3d72; assign y[491] = 16'hcebc;
	assign x[492] = 16'hb174; assign y[492] = 16'hfdf4;
	assign x[493] = 16'h1a30; assign y[493] = 16'h0a97;
	assign x[494] = 16'h8bcd; assign y[494] = 16'h118c;
	assign x[495] = 16'h8201; assign y[495] = 16'h945d;
	assign x[496] = 16'h6a08; assign y[496] = 16'hae39;
	assign x[497] = 16'hc5ab; assign y[497] = 16'h8053;
	assign x[498] = 16'h6afe; assign y[498] = 16'h3b63;
	assign x[499] = 16'ha8ac; assign y[499] = 16'h7c3c;
	assign x[500] = 16'hb4eb; assign y[500] = 16'h5339;
	assign x[501] = 16'h4e5d; assign y[501] = 16'ha94c;
	assign x[502] = 16'h04a7; assign y[502] = 16'h1a3e;
	assign x[503] = 16'h4ff5; assign y[503] = 16'hb06c;
	assign x[504] = 16'hb9f4; assign y[504] = 16'h9516;
	assign x[505] = 16'h963b; assign y[505] = 16'ha560;
	assign x[506] = 16'hfd5e; assign y[506] = 16'hceac;
	assign x[507] = 16'hdcac; assign y[507] = 16'h570e;
	assign x[508] = 16'h0084; assign y[508] = 16'h4811;
	assign x[509] = 16'h1652; assign y[509] = 16'he23f;
	assign x[510] = 16'h406f; assign y[510] = 16'haec4;
	assign x[511] = 16'h04c5; assign y[511] = 16'hf5f8;
	assign x[512] = 16'h83e4; assign y[512] = 16'h6014;
	assign x[513] = 16'h23f7; assign y[513] = 16'hd906;
	assign x[514] = 16'h8eb2; assign y[514] = 16'h5900;
	assign x[515] = 16'h56f7; assign y[515] = 16'h2067;
	assign x[516] = 16'h5096; assign y[516] = 16'h3858;
	assign x[517] = 16'hc4f7; assign y[517] = 16'hde88;
	assign x[518] = 16'h8811; assign y[518] = 16'h9f6f;
	assign x[519] = 16'h91e6; assign y[519] = 16'h06fb;
	assign x[520] = 16'hdb7f; assign y[520] = 16'h8f95;
	assign x[521] = 16'h8431; assign y[521] = 16'ha2c7;
	assign x[522] = 16'haf3d; assign y[522] = 16'h6146;
	assign x[523] = 16'hdd07; assign y[523] = 16'h488d;
	assign x[524] = 16'h0308; assign y[524] = 16'h4f87;
	assign x[525] = 16'hc4ae; assign y[525] = 16'hb8cd;
	assign x[526] = 16'heda2; assign y[526] = 16'h129e;
	assign x[527] = 16'hd2c2; assign y[527] = 16'h74e4;
	assign x[528] = 16'h0808; assign y[528] = 16'hb975;
	assign x[529] = 16'h5129; assign y[529] = 16'h6396;
	assign x[530] = 16'hb57d; assign y[530] = 16'hfe75;
	assign x[531] = 16'h09cc; assign y[531] = 16'h7f96;
	assign x[532] = 16'h7bf1; assign y[532] = 16'h8c87;
	assign x[533] = 16'h5eca; assign y[533] = 16'hd707;
	assign x[534] = 16'h27e5; assign y[534] = 16'he577;
	assign x[535] = 16'h7935; assign y[535] = 16'he639;
	assign x[536] = 16'h336a; assign y[536] = 16'h6066;
	assign x[537] = 16'h5437; assign y[537] = 16'he188;
	assign x[538] = 16'h2165; assign y[538] = 16'hda7e;
	assign x[539] = 16'hca1b; assign y[539] = 16'h8b30;
	assign x[540] = 16'h8160; assign y[540] = 16'hdfda;
	assign x[541] = 16'hb65b; assign y[541] = 16'ha7d0;
	assign x[542] = 16'h2e66; assign y[542] = 16'h9d31;
	assign x[543] = 16'h0f6d; assign y[543] = 16'hfc2b;
	assign x[544] = 16'h059d; assign y[544] = 16'h8049;
	assign x[545] = 16'h67d3; assign y[545] = 16'hcbb9;
	assign x[546] = 16'hc5f3; assign y[546] = 16'hdf08;
	assign x[547] = 16'hc74d; assign y[547] = 16'h13ab;
	assign x[548] = 16'hee3d; assign y[548] = 16'hb58b;
	assign x[549] = 16'h40ed; assign y[549] = 16'h8e83;
	assign x[550] = 16'ha7fe; assign y[550] = 16'h0c71;
	assign x[551] = 16'hcbd2; assign y[551] = 16'hf28c;
	assign x[552] = 16'h454b; assign y[552] = 16'h154a;
	assign x[553] = 16'h29b8; assign y[553] = 16'hb1e2;
	assign x[554] = 16'hb8d7; assign y[554] = 16'h024c;
	assign x[555] = 16'h2384; assign y[555] = 16'h61ad;
	assign x[556] = 16'h38bc; assign y[556] = 16'hf134;
	assign x[557] = 16'h1613; assign y[557] = 16'ha10a;
	assign x[558] = 16'h0cff; assign y[558] = 16'ha12d;
	assign x[559] = 16'hc909; assign y[559] = 16'h4023;
	assign x[560] = 16'h8cd7; assign y[560] = 16'hd015;
	assign x[561] = 16'h48c5; assign y[561] = 16'h4b83;
	assign x[562] = 16'hcef3; assign y[562] = 16'h9cb8;
	assign x[563] = 16'h1ea4; assign y[563] = 16'h5369;
	assign x[564] = 16'h4032; assign y[564] = 16'h4495;
	assign x[565] = 16'hf637; assign y[565] = 16'h17ea;
	assign x[566] = 16'h1641; assign y[566] = 16'hc647;
	assign x[567] = 16'h5c45; assign y[567] = 16'hb07c;
	assign x[568] = 16'h2a64; assign y[568] = 16'h2955;
	assign x[569] = 16'h594e; assign y[569] = 16'h87fa;
	assign x[570] = 16'h6738; assign y[570] = 16'h859d;
	assign x[571] = 16'ha7e7; assign y[571] = 16'h81fc;
	assign x[572] = 16'h84bb; assign y[572] = 16'he9b7;
	assign x[573] = 16'h4f76; assign y[573] = 16'he5cc;
	assign x[574] = 16'h4e3e; assign y[574] = 16'h13c3;
	assign x[575] = 16'h5a9b; assign y[575] = 16'h114d;
	assign x[576] = 16'ha1d5; assign y[576] = 16'h24ae;
	assign x[577] = 16'h62c2; assign y[577] = 16'he9c0;
	assign x[578] = 16'h7a39; assign y[578] = 16'head6;
	assign x[579] = 16'h519b; assign y[579] = 16'haad6;
	assign x[580] = 16'h450e; assign y[580] = 16'hf3f5;
	assign x[581] = 16'h1d44; assign y[581] = 16'h2a32;
	assign x[582] = 16'hafcf; assign y[582] = 16'h0142;
	assign x[583] = 16'h28f4; assign y[583] = 16'h353d;
	assign x[584] = 16'hdaff; assign y[584] = 16'hb463;
	assign x[585] = 16'he735; assign y[585] = 16'habee;
	assign x[586] = 16'hc191; assign y[586] = 16'hb95f;
	assign x[587] = 16'h3cd9; assign y[587] = 16'h45b0;
	assign x[588] = 16'ha23f; assign y[588] = 16'h0ba2;
	assign x[589] = 16'h5d7d; assign y[589] = 16'h400d;
	assign x[590] = 16'h09d4; assign y[590] = 16'hacff;
	assign x[591] = 16'h62fd; assign y[591] = 16'h1699;
	assign x[592] = 16'hd3e2; assign y[592] = 16'h1fc3;
	assign x[593] = 16'h9f5c; assign y[593] = 16'hc76e;
	assign x[594] = 16'h1abe; assign y[594] = 16'h5619;
	assign x[595] = 16'hb73c; assign y[595] = 16'h27a3;
	assign x[596] = 16'hd103; assign y[596] = 16'h1ba6;
	assign x[597] = 16'he1a4; assign y[597] = 16'hb5bf;
	assign x[598] = 16'h82fb; assign y[598] = 16'h9e96;
	assign x[599] = 16'he843; assign y[599] = 16'hd30f;
	assign x[600] = 16'h5c80; assign y[600] = 16'h0fb6;
	assign x[601] = 16'he84f; assign y[601] = 16'h873e;
	assign x[602] = 16'h6188; assign y[602] = 16'hc67b;
	assign x[603] = 16'h20d0; assign y[603] = 16'hb718;
	assign x[604] = 16'h314e; assign y[604] = 16'h3f29;
	assign x[605] = 16'h0d68; assign y[605] = 16'hb39a;
	assign x[606] = 16'h0aec; assign y[606] = 16'h5aab;
	assign x[607] = 16'hceba; assign y[607] = 16'h06fc;
	assign x[608] = 16'ha546; assign y[608] = 16'he9b7;
	assign x[609] = 16'hfdf7; assign y[609] = 16'hf3fc;
	assign x[610] = 16'h2930; assign y[610] = 16'h1a7b;
	assign x[611] = 16'hcdca; assign y[611] = 16'h8644;
	assign x[612] = 16'h0e3b; assign y[612] = 16'h3101;
	assign x[613] = 16'h2901; assign y[613] = 16'haacf;
	assign x[614] = 16'hb793; assign y[614] = 16'h326c;
	assign x[615] = 16'hf159; assign y[615] = 16'h10ee;
	assign x[616] = 16'h4efc; assign y[616] = 16'h92fc;
	assign x[617] = 16'h12d7; assign y[617] = 16'h005f;
	assign x[618] = 16'hc0dd; assign y[618] = 16'hace5;
	assign x[619] = 16'h5050; assign y[619] = 16'h4b34;
	assign x[620] = 16'h5234; assign y[620] = 16'h5967;
	assign x[621] = 16'h5165; assign y[621] = 16'h7c33;
	assign x[622] = 16'ha813; assign y[622] = 16'h0c35;
	assign x[623] = 16'hf740; assign y[623] = 16'hcbd4;
	assign x[624] = 16'h169d; assign y[624] = 16'h73ee;
	assign x[625] = 16'h7b07; assign y[625] = 16'h902a;
	assign x[626] = 16'ha83a; assign y[626] = 16'h570c;
	assign x[627] = 16'h79f3; assign y[627] = 16'hb444;
	assign x[628] = 16'h73bb; assign y[628] = 16'h53c6;
	assign x[629] = 16'hd76c; assign y[629] = 16'hed01;
	assign x[630] = 16'hba00; assign y[630] = 16'h46a7;
	assign x[631] = 16'hc5e4; assign y[631] = 16'h06e5;
	assign x[632] = 16'h5304; assign y[632] = 16'h02e2;
	assign x[633] = 16'hc7a1; assign y[633] = 16'h580b;
	assign x[634] = 16'h4c39; assign y[634] = 16'h09fd;
	assign x[635] = 16'h0ce2; assign y[635] = 16'ha58a;
	assign x[636] = 16'h01e4; assign y[636] = 16'h138c;
	assign x[637] = 16'h182b; assign y[637] = 16'h394b;
	assign x[638] = 16'h4b9e; assign y[638] = 16'h4e69;
	assign x[639] = 16'hc27e; assign y[639] = 16'h0d89;
	assign x[640] = 16'hd664; assign y[640] = 16'hdf5d;
	assign x[641] = 16'haa74; assign y[641] = 16'h7ef4;
	assign x[642] = 16'h4691; assign y[642] = 16'hba61;
	assign x[643] = 16'h6eee; assign y[643] = 16'hccff;
	assign x[644] = 16'h2566; assign y[644] = 16'h4274;
	assign x[645] = 16'hd0c5; assign y[645] = 16'hb380;
	assign x[646] = 16'h316f; assign y[646] = 16'hdcf2;
	assign x[647] = 16'hdf40; assign y[647] = 16'h7dc5;
	assign x[648] = 16'hf138; assign y[648] = 16'hc375;
	assign x[649] = 16'h7337; assign y[649] = 16'hca28;
	assign x[650] = 16'h7ae8; assign y[650] = 16'hf65d;
	assign x[651] = 16'hcb4b; assign y[651] = 16'h2356;
	assign x[652] = 16'h8136; assign y[652] = 16'h8d3f;
	assign x[653] = 16'hbe5c; assign y[653] = 16'h0b1f;
	assign x[654] = 16'hf2f8; assign y[654] = 16'h795a;
	assign x[655] = 16'h8d74; assign y[655] = 16'h14a2;
	assign x[656] = 16'ha4a4; assign y[656] = 16'hc813;
	assign x[657] = 16'h369c; assign y[657] = 16'h18f1;
	assign x[658] = 16'h49d5; assign y[658] = 16'hc8ec;
	assign x[659] = 16'h0db8; assign y[659] = 16'hd793;
	assign x[660] = 16'hc945; assign y[660] = 16'hddac;
	assign x[661] = 16'h35aa; assign y[661] = 16'hebdf;
	assign x[662] = 16'hec89; assign y[662] = 16'h52a0;
	assign x[663] = 16'h56d6; assign y[663] = 16'hae55;
	assign x[664] = 16'hf2df; assign y[664] = 16'hd27b;
	assign x[665] = 16'h5169; assign y[665] = 16'h9142;
	assign x[666] = 16'h399b; assign y[666] = 16'hbc8f;
	assign x[667] = 16'hb0da; assign y[667] = 16'h490f;
	assign x[668] = 16'hb71a; assign y[668] = 16'hf202;
	assign x[669] = 16'h1b99; assign y[669] = 16'h6431;
	assign x[670] = 16'h83e8; assign y[670] = 16'h5a92;
	assign x[671] = 16'ha63b; assign y[671] = 16'h9792;
	assign x[672] = 16'hc29e; assign y[672] = 16'h153a;
	assign x[673] = 16'h950c; assign y[673] = 16'hdcc7;
	assign x[674] = 16'h11de; assign y[674] = 16'hd233;
	assign x[675] = 16'h89c3; assign y[675] = 16'hc015;
	assign x[676] = 16'h6a95; assign y[676] = 16'hb199;
	assign x[677] = 16'h44b0; assign y[677] = 16'h43a9;
	assign x[678] = 16'h3879; assign y[678] = 16'hb6c3;
	assign x[679] = 16'h54de; assign y[679] = 16'h0ffc;
	assign x[680] = 16'hdc74; assign y[680] = 16'hcbfa;
	assign x[681] = 16'hed52; assign y[681] = 16'h26ff;
	assign x[682] = 16'h27d8; assign y[682] = 16'hd9d1;
	assign x[683] = 16'h46cf; assign y[683] = 16'h56a5;
	assign x[684] = 16'h4e51; assign y[684] = 16'h6a38;
	assign x[685] = 16'h5435; assign y[685] = 16'h74dd;
	assign x[686] = 16'h0f37; assign y[686] = 16'h4567;
	assign x[687] = 16'hfc70; assign y[687] = 16'hb6c5;
	assign x[688] = 16'h9379; assign y[688] = 16'hab9b;
	assign x[689] = 16'h3ca9; assign y[689] = 16'hd157;
	assign x[690] = 16'h8606; assign y[690] = 16'h510f;
	assign x[691] = 16'haf58; assign y[691] = 16'ha9e0;
	assign x[692] = 16'h4a06; assign y[692] = 16'hc095;
	assign x[693] = 16'h9c48; assign y[693] = 16'h7815;
	assign x[694] = 16'hc1d3; assign y[694] = 16'hb16b;
	assign x[695] = 16'hc7d0; assign y[695] = 16'hf14a;
	assign x[696] = 16'h9cc0; assign y[696] = 16'hd1f8;
	assign x[697] = 16'hd006; assign y[697] = 16'h3207;
	assign x[698] = 16'h4eda; assign y[698] = 16'h4b98;
	assign x[699] = 16'h0284; assign y[699] = 16'h36b0;
	assign x[700] = 16'h68eb; assign y[700] = 16'h38ed;
	assign x[701] = 16'h888a; assign y[701] = 16'h5657;
	assign x[702] = 16'hc070; assign y[702] = 16'h2bb6;
	assign x[703] = 16'h1271; assign y[703] = 16'h055e;
	assign x[704] = 16'h3b15; assign y[704] = 16'hb96d;
	assign x[705] = 16'hf61e; assign y[705] = 16'ha2ff;
	assign x[706] = 16'h375e; assign y[706] = 16'he7be;
	assign x[707] = 16'hbcf9; assign y[707] = 16'h81fd;
	assign x[708] = 16'hf91a; assign y[708] = 16'h751a;
	assign x[709] = 16'h516e; assign y[709] = 16'h27e6;
	assign x[710] = 16'h5604; assign y[710] = 16'h0d33;
	assign x[711] = 16'h5568; assign y[711] = 16'hd15b;
	assign x[712] = 16'h6a89; assign y[712] = 16'he059;
	assign x[713] = 16'hcf5e; assign y[713] = 16'h873b;
	assign x[714] = 16'h0ad6; assign y[714] = 16'h44be;
	assign x[715] = 16'hc6c4; assign y[715] = 16'h57b9;
	assign x[716] = 16'he1c5; assign y[716] = 16'h1b78;
	assign x[717] = 16'hc006; assign y[717] = 16'h2c70;
	assign x[718] = 16'hcf74; assign y[718] = 16'hab47;
	assign x[719] = 16'h7758; assign y[719] = 16'he93a;
	assign x[720] = 16'h1405; assign y[720] = 16'hf5bb;
	assign x[721] = 16'h341f; assign y[721] = 16'h8991;
	assign x[722] = 16'hfb05; assign y[722] = 16'hc9c6;
	assign x[723] = 16'hf202; assign y[723] = 16'h87d6;
	assign x[724] = 16'h5cae; assign y[724] = 16'h75a4;
	assign x[725] = 16'hba88; assign y[725] = 16'h51af;
	assign x[726] = 16'h9adb; assign y[726] = 16'h498b;
	assign x[727] = 16'he9f1; assign y[727] = 16'h233f;
	assign x[728] = 16'h2311; assign y[728] = 16'hf4cb;
	assign x[729] = 16'hc957; assign y[729] = 16'hd1e9;
	assign x[730] = 16'h2f3a; assign y[730] = 16'h87f3;
	assign x[731] = 16'hf6ee; assign y[731] = 16'h7594;
	assign x[732] = 16'h38c4; assign y[732] = 16'h97e8;
	assign x[733] = 16'h483a; assign y[733] = 16'hb80b;
	assign x[734] = 16'h3034; assign y[734] = 16'h46fa;
	assign x[735] = 16'h1d08; assign y[735] = 16'h460b;
	assign x[736] = 16'h65a2; assign y[736] = 16'h039c;
	assign x[737] = 16'h10ed; assign y[737] = 16'hcf07;
	assign x[738] = 16'hfb0e; assign y[738] = 16'h36ce;
	assign x[739] = 16'hf228; assign y[739] = 16'hb1ce;
	assign x[740] = 16'hafa3; assign y[740] = 16'h31ef;
	assign x[741] = 16'h02a2; assign y[741] = 16'h7bbe;
	assign x[742] = 16'h740b; assign y[742] = 16'hfed7;
	assign x[743] = 16'h9f7c; assign y[743] = 16'h8c85;
	assign x[744] = 16'h7300; assign y[744] = 16'h0497;
	assign x[745] = 16'hfdc3; assign y[745] = 16'hb5b0;
	assign x[746] = 16'hae86; assign y[746] = 16'h2eee;
	assign x[747] = 16'h27ae; assign y[747] = 16'h9c0a;
	assign x[748] = 16'hd836; assign y[748] = 16'h73d7;
	assign x[749] = 16'hbc28; assign y[749] = 16'hc327;
	assign x[750] = 16'h4a7b; assign y[750] = 16'h7698;
	assign x[751] = 16'h9367; assign y[751] = 16'h660c;
	assign x[752] = 16'hf655; assign y[752] = 16'hb7e4;
	assign x[753] = 16'h90d8; assign y[753] = 16'hc4c8;
	assign x[754] = 16'h423c; assign y[754] = 16'h3d29;
	assign x[755] = 16'hcd69; assign y[755] = 16'hb5ca;
	assign x[756] = 16'hf122; assign y[756] = 16'h7511;
	assign x[757] = 16'hbf74; assign y[757] = 16'hb7ae;
	assign x[758] = 16'hdd24; assign y[758] = 16'h8e08;
	assign x[759] = 16'hb7ea; assign y[759] = 16'hcd3f;
	assign x[760] = 16'h90f3; assign y[760] = 16'h35e8;
	assign x[761] = 16'hf59e; assign y[761] = 16'h952d;
	assign x[762] = 16'h3dc2; assign y[762] = 16'he458;
	assign x[763] = 16'h4efb; assign y[763] = 16'hb022;
	assign x[764] = 16'h7cb0; assign y[764] = 16'h5fb6;
	assign x[765] = 16'had1a; assign y[765] = 16'hffa4;
	assign x[766] = 16'h7517; assign y[766] = 16'h384e;
	assign x[767] = 16'hc48f; assign y[767] = 16'hc705;
	assign x[768] = 16'hedfc; assign y[768] = 16'hec6d;
	assign x[769] = 16'h70f9; assign y[769] = 16'hcc6f;
	assign x[770] = 16'h9f56; assign y[770] = 16'hf92d;
	assign x[771] = 16'h771e; assign y[771] = 16'ha109;
	assign x[772] = 16'h00d7; assign y[772] = 16'h2f0c;
	assign x[773] = 16'hf18b; assign y[773] = 16'ha260;
	assign x[774] = 16'hc9dd; assign y[774] = 16'h746a;
	assign x[775] = 16'hdcda; assign y[775] = 16'h18e5;
	assign x[776] = 16'h14b4; assign y[776] = 16'hd021;
	assign x[777] = 16'h2fdc; assign y[777] = 16'h86e4;
	assign x[778] = 16'h668d; assign y[778] = 16'ha753;
	assign x[779] = 16'h5b6d; assign y[779] = 16'h39e9;
	assign x[780] = 16'h5c94; assign y[780] = 16'hba72;
	assign x[781] = 16'h0e78; assign y[781] = 16'h77ab;
	assign x[782] = 16'h165f; assign y[782] = 16'h0424;
	assign x[783] = 16'hc3ed; assign y[783] = 16'h024e;
	assign x[784] = 16'h4262; assign y[784] = 16'h3ba4;
	assign x[785] = 16'h6613; assign y[785] = 16'h29c2;
	assign x[786] = 16'heea3; assign y[786] = 16'h6539;
	assign x[787] = 16'h00c3; assign y[787] = 16'hd495;
	assign x[788] = 16'h2230; assign y[788] = 16'h5ab1;
	assign x[789] = 16'h77f6; assign y[789] = 16'h7432;
	assign x[790] = 16'hd4b2; assign y[790] = 16'hc38c;
	assign x[791] = 16'hf309; assign y[791] = 16'h0030;
	assign x[792] = 16'hdf22; assign y[792] = 16'h6b92;
	assign x[793] = 16'hc332; assign y[793] = 16'h1517;
	assign x[794] = 16'h89e4; assign y[794] = 16'h0e9e;
	assign x[795] = 16'hb1b2; assign y[795] = 16'hbc24;
	assign x[796] = 16'hacb5; assign y[796] = 16'he867;
	assign x[797] = 16'h44cd; assign y[797] = 16'h2f21;
	assign x[798] = 16'h80e1; assign y[798] = 16'h34de;
	assign x[799] = 16'h34fc; assign y[799] = 16'h8bb5;
	assign x[800] = 16'h0c5a; assign y[800] = 16'h48a6;
	assign x[801] = 16'h4595; assign y[801] = 16'hc200;
	assign x[802] = 16'h6a07; assign y[802] = 16'ha39a;
	assign x[803] = 16'h673f; assign y[803] = 16'hd7a3;
	assign x[804] = 16'h3d9d; assign y[804] = 16'h3608;
	assign x[805] = 16'hf300; assign y[805] = 16'h3fc4;
	assign x[806] = 16'he537; assign y[806] = 16'hf089;
	assign x[807] = 16'h5b7b; assign y[807] = 16'he8e8;
	assign x[808] = 16'hadfc; assign y[808] = 16'h41fc;
	assign x[809] = 16'hd51a; assign y[809] = 16'h8245;
	assign x[810] = 16'hc124; assign y[810] = 16'h2837;
	assign x[811] = 16'habd2; assign y[811] = 16'h7795;
	assign x[812] = 16'he858; assign y[812] = 16'h7f37;
	assign x[813] = 16'hb3bc; assign y[813] = 16'hf60a;
	assign x[814] = 16'hd210; assign y[814] = 16'h0c3e;
	assign x[815] = 16'he4dd; assign y[815] = 16'h0313;
	assign x[816] = 16'hcf49; assign y[816] = 16'he464;
	assign x[817] = 16'h72ad; assign y[817] = 16'hdbe5;
	assign x[818] = 16'h7b6c; assign y[818] = 16'h81a5;
	assign x[819] = 16'hf457; assign y[819] = 16'hf33f;
	assign x[820] = 16'h4830; assign y[820] = 16'h74de;
	assign x[821] = 16'he1be; assign y[821] = 16'h9129;
	assign x[822] = 16'hb84e; assign y[822] = 16'hf8ed;
	assign x[823] = 16'h4c30; assign y[823] = 16'h2cd4;
	assign x[824] = 16'h600d; assign y[824] = 16'h998c;
	assign x[825] = 16'h3ed9; assign y[825] = 16'h1e34;
	assign x[826] = 16'h4f6a; assign y[826] = 16'haf84;
	assign x[827] = 16'h12c8; assign y[827] = 16'hab3b;
	assign x[828] = 16'h521a; assign y[828] = 16'hefec;
	assign x[829] = 16'hc7d5; assign y[829] = 16'h6011;
	assign x[830] = 16'hd2ac; assign y[830] = 16'hfe00;
	assign x[831] = 16'h6254; assign y[831] = 16'h55c4;
	assign x[832] = 16'hc823; assign y[832] = 16'h1821;
	assign x[833] = 16'had8c; assign y[833] = 16'h6012;
	assign x[834] = 16'ha7f6; assign y[834] = 16'h5dcc;
	assign x[835] = 16'hde3a; assign y[835] = 16'h4de6;
	assign x[836] = 16'hfca4; assign y[836] = 16'h6d3f;
	assign x[837] = 16'he1fc; assign y[837] = 16'h10d9;
	assign x[838] = 16'h7c66; assign y[838] = 16'hf9bb;
	assign x[839] = 16'ha2a7; assign y[839] = 16'h648d;
	assign x[840] = 16'h0043; assign y[840] = 16'h164b;
	assign x[841] = 16'h1fe1; assign y[841] = 16'h44b1;
	assign x[842] = 16'h7c56; assign y[842] = 16'he2ed;
	assign x[843] = 16'h72af; assign y[843] = 16'h37d5;
	assign x[844] = 16'hd9de; assign y[844] = 16'h92a2;
	assign x[845] = 16'had21; assign y[845] = 16'hfca2;
	assign x[846] = 16'h6260; assign y[846] = 16'h5390;
	assign x[847] = 16'hbeca; assign y[847] = 16'hb68b;
	assign x[848] = 16'he054; assign y[848] = 16'hc819;
	assign x[849] = 16'he0b7; assign y[849] = 16'ha292;
	assign x[850] = 16'hefe8; assign y[850] = 16'h2278;
	assign x[851] = 16'h4b0d; assign y[851] = 16'h7086;
	assign x[852] = 16'h3a02; assign y[852] = 16'h4fc1;
	assign x[853] = 16'hc9c1; assign y[853] = 16'hed81;
	assign x[854] = 16'h6b87; assign y[854] = 16'hbc5a;
	assign x[855] = 16'h17dc; assign y[855] = 16'h0ae4;
	assign x[856] = 16'hcff1; assign y[856] = 16'h6a26;
	assign x[857] = 16'h2cd5; assign y[857] = 16'hd31d;
	assign x[858] = 16'hd2a2; assign y[858] = 16'h6bc2;
	assign x[859] = 16'h021e; assign y[859] = 16'h45d3;
	assign x[860] = 16'hfabb; assign y[860] = 16'h9e04;
	assign x[861] = 16'hc2a2; assign y[861] = 16'h21d0;
	assign x[862] = 16'h2814; assign y[862] = 16'hfc48;
	assign x[863] = 16'h07d4; assign y[863] = 16'h686c;
	assign x[864] = 16'hd6b4; assign y[864] = 16'hb853;
	assign x[865] = 16'h9fc9; assign y[865] = 16'h2adc;
	assign x[866] = 16'h0be5; assign y[866] = 16'h7a6e;
	assign x[867] = 16'h0e47; assign y[867] = 16'hbc2a;
	assign x[868] = 16'h4e87; assign y[868] = 16'hee77;
	assign x[869] = 16'h844c; assign y[869] = 16'h386a;
	assign x[870] = 16'he4f1; assign y[870] = 16'h8e91;
	assign x[871] = 16'h7066; assign y[871] = 16'hc3f3;
	assign x[872] = 16'hc4a3; assign y[872] = 16'hadf6;
	assign x[873] = 16'h74e4; assign y[873] = 16'h871b;
	assign x[874] = 16'h2d8e; assign y[874] = 16'h1688;
	assign x[875] = 16'h4f40; assign y[875] = 16'ha18d;
	assign x[876] = 16'hf857; assign y[876] = 16'h2068;
	assign x[877] = 16'hf579; assign y[877] = 16'hde90;
	assign x[878] = 16'ha38d; assign y[878] = 16'hc564;
	assign x[879] = 16'h0c6f; assign y[879] = 16'h3bb2;
	assign x[880] = 16'hde55; assign y[880] = 16'h4464;
	assign x[881] = 16'h4892; assign y[881] = 16'h0fef;
	assign x[882] = 16'h3ce1; assign y[882] = 16'hdc0a;
	assign x[883] = 16'h7eea; assign y[883] = 16'h1046;
	assign x[884] = 16'h8b42; assign y[884] = 16'h8740;
	assign x[885] = 16'hc4c2; assign y[885] = 16'h3b19;
	assign x[886] = 16'hb009; assign y[886] = 16'h9550;
	assign x[887] = 16'hbf5a; assign y[887] = 16'h610b;
	assign x[888] = 16'h1e84; assign y[888] = 16'had70;
	assign x[889] = 16'h0724; assign y[889] = 16'h52a6;
	assign x[890] = 16'hfdac; assign y[890] = 16'h0b3d;
	assign x[891] = 16'h8405; assign y[891] = 16'ha9c4;
	assign x[892] = 16'h467c; assign y[892] = 16'hb026;
	assign x[893] = 16'h32da; assign y[893] = 16'hd5d6;
	assign x[894] = 16'h22a4; assign y[894] = 16'h80c7;
	assign x[895] = 16'h3558; assign y[895] = 16'h2671;
	assign x[896] = 16'h41ab; assign y[896] = 16'hf875;
	assign x[897] = 16'h11be; assign y[897] = 16'h7260;
	assign x[898] = 16'hb1d4; assign y[898] = 16'h3191;
	assign x[899] = 16'h6f16; assign y[899] = 16'h5ab8;
	assign x[900] = 16'h75d6; assign y[900] = 16'hcc4e;
	assign x[901] = 16'h671e; assign y[901] = 16'he0c2;
	assign x[902] = 16'hb263; assign y[902] = 16'h50e0;
	assign x[903] = 16'h89d1; assign y[903] = 16'hb273;
	assign x[904] = 16'h66ce; assign y[904] = 16'h6ea0;
	assign x[905] = 16'hee74; assign y[905] = 16'ha0a1;
	assign x[906] = 16'h41c6; assign y[906] = 16'h8dbb;
	assign x[907] = 16'h003b; assign y[907] = 16'h2aa3;
	assign x[908] = 16'ha7fa; assign y[908] = 16'h9de1;
	assign x[909] = 16'ha583; assign y[909] = 16'h11f9;
	assign x[910] = 16'h2b4c; assign y[910] = 16'h073a;
	assign x[911] = 16'h95b6; assign y[911] = 16'h3ab4;
	assign x[912] = 16'h553d; assign y[912] = 16'h8cf4;
	assign x[913] = 16'h671f; assign y[913] = 16'hb154;
	assign x[914] = 16'he5ef; assign y[914] = 16'h2d85;
	assign x[915] = 16'hd448; assign y[915] = 16'hd17f;
	assign x[916] = 16'h3ed3; assign y[916] = 16'h2926;
	assign x[917] = 16'hed08; assign y[917] = 16'ha5f4;
	assign x[918] = 16'h5928; assign y[918] = 16'h97d7;
	assign x[919] = 16'h7b69; assign y[919] = 16'hdfb8;
	assign x[920] = 16'h92ce; assign y[920] = 16'h100c;
	assign x[921] = 16'h0bba; assign y[921] = 16'h0435;
	assign x[922] = 16'h89e0; assign y[922] = 16'h2700;
	assign x[923] = 16'ha050; assign y[923] = 16'ha243;
	assign x[924] = 16'h932a; assign y[924] = 16'h18cc;
	assign x[925] = 16'h7f64; assign y[925] = 16'h47b0;
	assign x[926] = 16'h84e6; assign y[926] = 16'h1cb7;
	assign x[927] = 16'hc6f8; assign y[927] = 16'hd652;
	assign x[928] = 16'h8fce; assign y[928] = 16'h736c;
	assign x[929] = 16'h81c6; assign y[929] = 16'ha020;
	assign x[930] = 16'hfa9f; assign y[930] = 16'he5ca;
	assign x[931] = 16'h3eea; assign y[931] = 16'hd8e9;
	assign x[932] = 16'hbfba; assign y[932] = 16'h56cd;
	assign x[933] = 16'h1a41; assign y[933] = 16'h7647;
	assign x[934] = 16'hf463; assign y[934] = 16'hc474;
	assign x[935] = 16'h0fab; assign y[935] = 16'h7a1b;
	assign x[936] = 16'h2986; assign y[936] = 16'h9dd9;
	assign x[937] = 16'h3264; assign y[937] = 16'h5d80;
	assign x[938] = 16'h41e2; assign y[938] = 16'he016;
	assign x[939] = 16'h07c7; assign y[939] = 16'hb96e;
	assign x[940] = 16'hd3eb; assign y[940] = 16'h3fc6;
	assign x[941] = 16'h7e39; assign y[941] = 16'hffea;
	assign x[942] = 16'h9039; assign y[942] = 16'h897f;
	assign x[943] = 16'hcef5; assign y[943] = 16'hdcee;
	assign x[944] = 16'hf102; assign y[944] = 16'h1de0;
	assign x[945] = 16'h5416; assign y[945] = 16'hb6f0;
	assign x[946] = 16'h67a9; assign y[946] = 16'h7f99;
	assign x[947] = 16'h4d63; assign y[947] = 16'h714f;
	assign x[948] = 16'h9a07; assign y[948] = 16'h4a64;
	assign x[949] = 16'h5f60; assign y[949] = 16'h8034;
	assign x[950] = 16'h0df3; assign y[950] = 16'h5ccc;
	assign x[951] = 16'h771b; assign y[951] = 16'hd5b1;
	assign x[952] = 16'h504d; assign y[952] = 16'h7c98;
	assign x[953] = 16'h41f4; assign y[953] = 16'h5604;
	assign x[954] = 16'h7ef3; assign y[954] = 16'h9949;
	assign x[955] = 16'h0ac5; assign y[955] = 16'hebf8;
	assign x[956] = 16'h664a; assign y[956] = 16'h1fee;
	assign x[957] = 16'hd2f7; assign y[957] = 16'h55eb;
	assign x[958] = 16'hc314; assign y[958] = 16'hc69b;
	assign x[959] = 16'h6ccb; assign y[959] = 16'hc505;
	assign x[960] = 16'hfc82; assign y[960] = 16'h34c1;
	assign x[961] = 16'h40e8; assign y[961] = 16'h2c03;
	assign x[962] = 16'h05f7; assign y[962] = 16'h29da;
	assign x[963] = 16'h0566; assign y[963] = 16'h7c6e;
	assign x[964] = 16'hcaaf; assign y[964] = 16'he698;
	assign x[965] = 16'h8d34; assign y[965] = 16'hd32c;
	assign x[966] = 16'hb0ca; assign y[966] = 16'hcae7;
	assign x[967] = 16'h8439; assign y[967] = 16'h273c;
	assign x[968] = 16'h50c0; assign y[968] = 16'h7c3f;
	assign x[969] = 16'h6b77; assign y[969] = 16'h1737;
	assign x[970] = 16'h1b79; assign y[970] = 16'h2252;
	assign x[971] = 16'he47b; assign y[971] = 16'h7f7b;
	assign x[972] = 16'he6b6; assign y[972] = 16'h44db;
	assign x[973] = 16'h940c; assign y[973] = 16'h06e8;
	assign x[974] = 16'h4ba4; assign y[974] = 16'hb3d0;
	assign x[975] = 16'hb749; assign y[975] = 16'hbbea;
	assign x[976] = 16'h983e; assign y[976] = 16'h81cb;
	assign x[977] = 16'h4469; assign y[977] = 16'h0b85;
	assign x[978] = 16'hf57a; assign y[978] = 16'h6632;
	assign x[979] = 16'hcb37; assign y[979] = 16'hadc2;
	assign x[980] = 16'hf272; assign y[980] = 16'h9a53;
	assign x[981] = 16'he178; assign y[981] = 16'h4755;
	assign x[982] = 16'hf36d; assign y[982] = 16'h9780;
	assign x[983] = 16'ha9eb; assign y[983] = 16'hb2b0;
	assign x[984] = 16'hc2eb; assign y[984] = 16'hcaae;
	assign x[985] = 16'hcd73; assign y[985] = 16'h9886;
	assign x[986] = 16'h7871; assign y[986] = 16'h60ab;
	assign x[987] = 16'hdcd6; assign y[987] = 16'h6eca;
	assign x[988] = 16'h87c2; assign y[988] = 16'h55b6;
	assign x[989] = 16'h47d0; assign y[989] = 16'hf3a3;
	assign x[990] = 16'haef5; assign y[990] = 16'h8498;
	assign x[991] = 16'hdde9; assign y[991] = 16'h9a72;
	assign x[992] = 16'he994; assign y[992] = 16'h1ab4;
	assign x[993] = 16'h637e; assign y[993] = 16'h8394;
	assign x[994] = 16'heaea; assign y[994] = 16'h2336;
	assign x[995] = 16'h095b; assign y[995] = 16'h670b;
	assign x[996] = 16'h34d8; assign y[996] = 16'h8340;
	assign x[997] = 16'h0089; assign y[997] = 16'h6ee3;
	assign x[998] = 16'h5eb8; assign y[998] = 16'h58e0;
	assign x[999] = 16'hb883; assign y[999] = 16'h890c;

	initial begin
		$display("test: testmul");
		for (i = 0; i < $size(x); i = i + 1) begin
			xin = x[i];
			yin = y[i];
			zmul = xin * yin;
			#10;
			if (zmul != z)
				$display("xin=0x%4H yin=0x%4H got=%8H expected=%8H", xin, yin, z, zmul);
		end
		$finish;
	end
endmodule
