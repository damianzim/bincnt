// vim: ts=4 sts=0 sw=0 noet
`default_nettype none
`timescale 1ns / 1ns

module ha (
	input wire [1:0] x,
	output wire [1:0] y
);
	assign y = {x[0]&x[1], x[0]^x[1]};
endmodule

module fa (
	input wire [2:0] x,
	output wire [1:0] y
);
	assign y = {(x[0]&x[1])|((x[0]^x[1])&x[2]), (x[0]^x[1])^x[2]};
endmodule

module multiplier16b (
	input wire [15:0] x, y,
	output wire [31:0] z
);
	wire [15:0][15:0] l1;

	assign l1[0] = y[0] == 0 ? '0 : x;
	assign l1[1] = y[1] == 0 ? '0 : x;
	assign l1[2] = y[2] == 0 ? '0 : x;
	assign l1[3] = y[3] == 0 ? '0 : x;
	assign l1[4] = y[4] == 0 ? '0 : x;
	assign l1[5] = y[5] == 0 ? '0 : x;
	assign l1[6] = y[6] == 0 ? '0 : x;
	assign l1[7] = y[7] == 0 ? '0 : x;
	assign l1[8] = y[8] == 0 ? '0 : x;
	assign l1[9] = y[9] == 0 ? '0 : x;
	assign l1[10] = y[10] == 0 ? '0 : x;
	assign l1[11] = y[11] == 0 ? '0 : x;
	assign l1[12] = y[12] == 0 ? '0 : x;
	assign l1[13] = y[13] == 0 ? '0 : x;
	assign l1[14] = y[14] == 0 ? '0 : x;
	assign l1[15] = y[15] == 0 ? '0 : x;

	wire l2p0 = l1[0][0];
	wire l2p1;
	wire [1:0] l2p2;
	wire [1:0] l2p3;
	wire [1:0] l2p4;
	wire [2:0] l2p5;
	wire [2:0] l2p6;
	wire [3:0] l2p7;
	wire [4:0] l2p8;
	wire [3:0] l2p9;
	wire [4:0] l2p10;
	wire [4:0] l2p11;
	wire [5:0] l2p12;
	wire [5:0] l2p13;
	wire [6:0] l2p14;
	wire [6:0] l2p15;
	wire [6:0] l2p16;
	wire [6:0] l2p17;
	wire [5:0] l2p18;
	wire [5:0] l2p19;
	wire [5:0] l2p20;
	wire [5:0] l2p21;
	wire [6:0] l2p22;
	wire [3:0] l2p23;
	wire [2:0] l2p24;
	wire [2:0] l2p25;
	wire [2:0] l2p26;
	wire [2:0] l2p27;
	wire [2:0] l2p28;
	wire [2:0] l2p29;
	wire [1:0] l2p30;

	// ===== BEGIN L1 =====
	ha hal1p1 (.x ({l1[0][1], l1[1][0]}), .y ({l2p2[0], l2p1})); // R: l2p2[0:0], l2p1
	fa fal1p2 (.x ({l1[0][2], l1[1][1], l1[2][0]}), .y ({l2p3[0], l2p2[1]})); // R: l2p3[0], l2p2[1:0]
	counter7b3 cnt7bl1p3 (
		.x ({l1[0][3], l1[1][2], l1[2][1], l1[3][0], 3'b000}),
		.y ({l2p5[0], l2p4[0], l2p3[1]})
	); // R: l2p5[0], l2p4[0], l2p3[1:0]
	counter7b3 cnt7bl1p4 (
		.x ({l1[0][4], l1[1][3], l1[2][2], l1[3][1], l1[4][0], 2'b00}),
		.y ({l2p6[0], l2p5[1], l2p4[1]})
	); // R:l2p6[0], l2p5[1:0], l2p4[1:0]
	counter7b3 cnt7bl1p5 (
		.x ({l1[0][5], l1[1][4], l1[2][3], l1[3][2], l1[4][1], l1[5][0], 1'b0}),
		.y ({l2p7[0], l2p6[1], l2p5[2]})
	); // R: l2p7[0], l2p6[1:0], l2p5[2:0]
	counter7b3 cnt7bl1p6 (
		.x ({l1[0][6], l1[1][5], l1[2][4], l1[3][3], l1[4][2], l1[5][1], l1[6][0]}),
		.y ({l2p8[0], l2p7[1], l2p6[2]})
	); // R:l2p8[0], l2p7[1:0], l2p6[2:0]
	counter7b3 cnt7bl1p7 (
		.x ({l1[0][7], l1[1][6], l1[2][5], l1[3][4], l1[4][3], l1[5][2], l1[6][1]}),
		.y ({l2p9[0], l2p8[1], l2p7[2]})
	); // R: l2p9[0], l2p8[1:0], l2p7[2:0]
	assign l2p7[3] = l1[7][0]; // R: l2p7[3:0]
	counter7b3 cnt7bl1p8 (
		.x ({l1[0][8], l1[1][7], l1[2][6], l1[3][5], l1[4][4], l1[5][3], l1[6][2]}),
		.y ({l2p10[0], l2p9[1], l2p8[2]})
	); // R: l2p10[0], l2p9[1:0], l2p8[2:0]
	assign l2p8[4:3] = {l1[7][1], l1[8][0]};
	counter7b3 cnt7bl1p9 (
		.x ({l1[0][9], l1[1][8], l1[2][7], l1[3][6], l1[4][5], l1[5][4], l1[6][3]}),
		.y ({l2p11[0], l2p10[1], l2p9[2]})
	); // R: l2p11[0], l2p10[1:0], l2p9[2:0]
	fa fal1p9 (
		.x ({l1[7][2], l1[8][1], l1[9][0]}),
		.y ({l2p10[2], l2p9[3]})
	); // R: l2p10[2:0], l2p9[3:0]
	counter7b3 cnt7bl1p10_0 (
		.x ({l1[0][10], l1[1][9], l1[2][8], l1[3][7], l1[4][6], l1[5][5], l1[6][4]}),
		.y ({l2p12[0], l2p11[1], l2p10[3]})
	); // R: l2p12[0], l2p11[1:0], l2p10[3:0]
	counter7b3 cnt7bl1p10_1 (
		.x ({l1[7][3], l1[8][2], l1[9][1], l1[10][0], 3'b000}),
		.y ({l2p12[1], l2p11[2], l2p10[4]})
	); // R: l2p12[1:0], l2p11[2:0], l2p10[4:0]
	counter7b3 cnt7bl1p11_0 (
		.x ({l1[0][11], l1[1][10], l1[2][9], l1[3][8], l1[4][7], l1[5][6], l1[6][5]}),
		.y ({l2p13[0], l2p12[2], l2p11[3]})
	); // R: l2p13[0], l2p12[2:0], l2p11[3:0]
	counter7b3 cnt7bl1p11_1 (
		.x ({l1[7][4], l1[8][3], l1[9][2], l1[10][1], l1[11][0], 2'b00}),
		.y ({l2p13[1], l2p12[3], l2p11[4]})
	); // R: l2p13[1:0], l2p12[3:0], l2p11[4:0]
	counter7b3 cnt7bl1p12_0 (
		.x ({l1[0][12], l1[1][11], l1[2][10], l1[3][9], l1[4][8], l1[5][7], l1[6][6]}),
		.y ({l2p14[0], l2p11[2], l2p12[4]})
	); // R: l2p14[0], l2p13[2:0], l2p12[4:0]
	counter7b3 cnt7bl1p12_1 (
		.x ({l1[7][5], l1[8][4], l1[9][3], l1[10][2], l1[11][1], l1[12][0], 1'b0}),
		.y ({l2p14[1], l2p13[3], l2p12[5]})
	); // R: l2p14[1:0], l2p13[3:0], l2p12[5:0]
	counter7b3 cnt7bl1p13_0 (
		.x ({l1[0][13], l1[1][12], l1[2][11], l1[3][10], l1[4][9], l1[5][8], l1[6][7]}),
		.y ({l2p15[0], l2p14[2], l2p13[4]})
	); // R: l2p15[0], l2p14[2:0], l2p13[4:0]
	counter7b3 cnt7bl1p13_1 (
		.x ({l1[7][6], l1[8][5], l1[9][4], l1[10][3], l1[11][2], l1[12][1], l1[13][0]}),
		.y ({l2p15[1], l2p14[3], l2p13[5]})
	); // R: l2p15[1:0], l2p14[3:0], l2p13[5:0]
	counter7b3 cnt7bl1p14_0 (
		.x ({l1[0][14], l1[1][13], l1[2][12], l1[3][11], l1[4][10], l1[5][9], l1[6][8]}),
		.y ({l2p16[0], l2p15[2], l2p14[4]})
	); // R: l2p16[0], l2p15[2:0], l2p14[4:0]
	counter7b3 cnt7bl1p14_1 (
		.x ({l1[7][7], l1[8][6], l1[9][5], l1[10][4], l1[11][3], l1[12][2], l1[13][1]}),
		.y ({l2p16[1], l2p15[3], l2p14[5]})
	); // R: l2p16[1:0], l2p15[3:0], l2p14[5:0]
	assign l2p14[6] = l1[14][0];
	counter7b3 cnt7bl1p15_0 (
		.x ({l1[0][15], l1[1][14], l1[2][13], l1[3][12], l1[4][11], l1[5][10], l1[6][9]}),
		.y ({l2p17[0], l2p16[2], l2p15[4]})
	); // R: l2p17[0], l2p16[2:0], l2p15[4:0]
	counter7b3 cnt7bl1p15_1 (
		.x ({l1[7][8], l1[8][7], l1[9][6], l1[10][5], l1[11][4], l1[12][3], l1[13][2]}),
		.y ({l2p17[1], l2p16[3], l2p15[5]})
	); // R: l2p17[1:0], l2p16[3:0], l2p15[5:0]
	counter7b3 cnt7bl1p15_2 (
		.x ({l1[14][1], l1[15][0], l1[15][1], l1[15][1], 3'b000}), // l1[15][1] is repeated, beacause it has weight x2
		.y ({l2p17[2], l2p16[4], l2p15[6]})
	); // R: l2p17[2:0], l2p16[4:0], l2p15[6:0]
	counter7b3 cnt7bl1p16_0 (
		.x ({l1[1][15], l1[2][14], l1[3][13], l1[4][12], l1[5][11], l1[6][10], l1[7][9]}),
		.y ({l2p18[0], l2p17[3], l2p16[5]})
	); // R: l2p18[0], l2p17[3:0], l2p16[5:0]
	counter7b3 cnt7bl1p16_1 (
		.x ({l1[8][8], l1[9][7], l1[10][6], l1[11][5], l1[12][4], l1[13][3], l1[14][2]}),
		.y ({l2p18[1], l2p17[4], l2p16[6]})
	); // R: l2p18[1:0], l2p17[4:0], l2p16[6:0]
	counter7b3 cnt7bl1p17_0 (
		.x ({l1[2][15], l1[3][14], l1[4][13], l1[5][12], l1[6][11], l1[7][10], l1[8][9]}),
		.y ({l2p19[0], l2p18[2], l2p17[5]})
	); // R: l2p19[0], l2p18[2:0], l2p17[5:0]
	counter7b3 cnt7bl1p17_1 (
		.x ({l1[9][8], l1[10][7], l1[11][6], l1[12][5], l1[13][4], l1[14][3], l1[15][3]}),
		.y ({l2p19[1], l2p18[3], l2p17[6]})
	); // R: l2p19[1:0], l2p18[3:0], l2p17[6:0]
	counter7b3 cnt7bl1p18_0 (
		.x ({l1[3][15], l1[4][14], l1[5][13], l1[6][12], l1[7][11], l1[8][10], l1[9][9]}),
		.y ({l2p20[0], l2p19[2], l2p18[4]})
	); // R: l2p20[0], l2p19[2:0], l2p18[4:0]
	counter7b3 cnt7bl1p18_1 (
		.x ({l1[10][8], l1[11][7], l1[12][6], l1[13][5], l1[14][4], l1[15][3], 1'b0}),
		.y ({l2p20[1], l2p19[3], l2p18[5]})
	); // R: l2p20[1:0], l2p19[3:0], l2p18[5:0]
	counter7b3 cnt7bl1p19_0 (
		.x ({l1[4][15], l1[5][14], l1[6][13], l1[7][12], l1[8][11], l1[9][10], l1[10][9]}),
		.y ({l2p21[0], l2p20[2], l2p19[4]})
	); // R: l2p21[0], l2p20[2:0], l2p19[4:0]
	counter7b3 cnt7bl1p19_1 (
		.x ({l1[11][8], l1[12][7], l1[13][6], l1[14][5], l1[15][4], 2'b00}),
		.y ({l2p21[1], l2p20[3], l2p19[5]})
	); // R: l2p21[1:0], l2p20[3:0], l2p19[5:0]
	counter7b3 cnt7bl1p20_0 (
		.x ({l1[5][15], l1[6][14], l1[7][13], l1[8][12], l1[9][11], l1[10][10], l1[11][9]}),
		.y ({l2p22[0], l2p21[2], l2p20[4]})
	); // R: l2p22[0], l2p21[2:0], l2p20[4:0]
	counter7b3 cnt7bl1p20_1 (
		.x ({l1[12][8], l1[13][7], l1[14][6], l1[15][5], 3'b000}),
		.y ({l2p22[1], l2p21[3], l2p20[5]})
	); // R: l2p22[1:0], l2p21[3:0], l2p20[5:0]
	counter7b3 cnt7bl1p21 (
		.x ({l1[6][15], l1[7][14], l1[8][13], l1[9][12], l1[10][11], l1[11][10], l1[12][9]}),
		.y ({l2p23[0], l2p22[2], l2p21[4]})
	); // R: l2p23[0], l2p22[2:0], l2p21[4:0]
	fa fal1p21 (
		.x ({l1[13][8], l1[14][7], l1[15][6]}),
		.y ({l2p22[3], l2p21[5]})
	); // R: l2p22[3:0], l2p21[5:0]
	counter7b3 cnt7bl1p22 (
		.x ({l1[7][15], l1[8][14], l1[9][13], l1[10][12], l1[11][11], l1[12][10], l1[13][9]}),
		.y ({l2p24[0], l2p23[1], l2p22[4]})
	); // R: l2p24[0], l2p23[1:0], l2p22[4:0]
	assign l2p22[6:5] = {l1[14][8], l1[15][7]}; // R: l2p22[6:0]
	counter7b3 cnt7bl1p23 (
		.x ({l1[8][15], l1[9][14], l1[10][13], l1[11][12], l1[12][11], l1[13][10], l1[14][9]}),
		.y ({l2p25[0], l2p24[1], l2p23[2]})
	); // R: l2p25[0], l2p24[1:0], l2p23[2:0]
	assign l2p23[3] = l1[15][8]; // R: l2p23[3:0]
	counter7b3 cnt7bl1p24 (
		.x ({l1[9][15], l1[10][14], l1[11][13], l1[12][12], l1[13][11], l1[14][10], l1[15][9]}),
		.y ({l2p26[0], l2p25[1], l2p24[2]})
	); // R: l2p26[0], l2p25[1:0], l2p24[2:0]
	counter7b3 cnt7bl1p25 (
		.x ({l1[10][15], l1[11][14], l1[12][13], l1[13][12], l1[14][11], l1[15][10], 1'b0}),
		.y ({l2p27[0], l2p26[1], l2p25[2]})
	); // R: l2p27[0], l2p26[1:0], l2p25[2:0]
	counter7b3 cnt7bl1p26 (
		.x ({l1[11][15], l1[12][14], l1[13][13], l1[14][12], l1[15][11], 2'b00}),
		.y ({l2p28[0], l2p27[1], l2p26[2]})
	); // R: l2p28[0], l2p27[1:0], l2p26[2:0]
	counter7b3 cnt7bl1p27 (
		.x ({l1[12][15], l1[13][14], l1[14][13], l1[15][12]}),
		.y ({l2p29[0], l2p28[1], l2p27[2]})
	); // R: l2p29[0], l2p28[1:0], l2p27[2:0]
	fa fal1p28 (
		.x ({l1[13][15], l1[14][14], l1[15][13]}),
		.y ({l2p29[1], l2p28[2]})
	); // R: l2p29[1:0], l2p28[2:0]
	ha hal1p29 (
		.x ({l1[14][15], l1[15][14]}),
		.y ({l2p30[0], l2p29[2]})
	); // R: l2p30[0], l2p29[2:0]
	assign l2p30[1] = l1[15][15];
	// ===== END L1 =====

	//assign z[15:0] = x;
	//assign z[31:16] = y;
endmodule
